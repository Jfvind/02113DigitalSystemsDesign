module Memory(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_1(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_2(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_2.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_3(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_3.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_4(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_4.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_5(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_5.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_6(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_6.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_7(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_7.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_8(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_8.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_9(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_9.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_10(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_10.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_11(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_11.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_12(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_12.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_13(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_13.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_14(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_14.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_15(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_15.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_16(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_16.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_17(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_17.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_18(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_18.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_19(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_19.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_20(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_20.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_21(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_21.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_22(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_22.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_23(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_23.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_24(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_24.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_25(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_25.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_26(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_26.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_27(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_27.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_28(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_28.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_29(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_29.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_30(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_30.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_31(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_31.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_32(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_32.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_33(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_33.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_34(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_34.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_35(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_35.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_36(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_36.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_37(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_37.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_38(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_38.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_39(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_39.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_40(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_40.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_41(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_41.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_42(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_42.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_43(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_43.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_44(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_44.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_45(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_45.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_46(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_46.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_47(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_47.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_48(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_48.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_49(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_49.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_50(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_50.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_51(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_51.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_52(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_52.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_53(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_53.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_54(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_54.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_55(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_55.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_56(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_56.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_57(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_57.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_58(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_58.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_59(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_59.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_60(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_60.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_61(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_61.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_62(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_62.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_63(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_63.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_64(
  input         clock,
  input  [10:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [5:0]  io_dataRead, // @[\\src\\main\\scala\\Memory.scala 48:14]
  input         io_writeEnable, // @[\\src\\main\\scala\\Memory.scala 48:14]
  input  [5:0]  io_dataWrite // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [10:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [5:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [5:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 57:26]
  RamSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(6)) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 57:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 63:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 58:21]
  assign ramsSpWf_we = io_writeEnable; // @[\\src\\main\\scala\\Memory.scala 59:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 60:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 61:22]
  assign ramsSpWf_di = io_dataWrite; // @[\\src\\main\\scala\\Memory.scala 62:20]
endmodule
module Memory_66(
  input         clock,
  input  [10:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [5:0]  io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [10:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [5:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [5:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(6), .LOAD_FILE("memory_init/backbuffer_init.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 6'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_67(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_68(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_69(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_2.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_70(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_3.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_71(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_4.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_72(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_5.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_73(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_6.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_74(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_7.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_75(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_8.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_76(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_9.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_77(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_10.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_78(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_11.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_79(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_12.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_80(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_13.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_81(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_14.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_82(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_15.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_83(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_16.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_84(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_17.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_85(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_18.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_86(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_19.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_87(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_20.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_88(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_21.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_89(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_22.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_90(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_23.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_91(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_24.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_92(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_25.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_93(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_26.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_94(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_27.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_95(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_28.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_96(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_29.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_97(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_30.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_98(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_31.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_99(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_32.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_100(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_33.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_101(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_34.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_102(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_35.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_103(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_36.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_104(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_37.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_105(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_38.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_106(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_39.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_107(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_40.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_108(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_41.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_109(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_42.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_110(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_43.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_111(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_44.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_112(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_45.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_113(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_46.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_114(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_47.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_115(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_48.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_116(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_49.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_117(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_50.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_118(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_51.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_119(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_52.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_120(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_53.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_121(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_54.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_122(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_55.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_123(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_56.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_124(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_57.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_125(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_58.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_126(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_59.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_127(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_60.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_128(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_61.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_129(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_62.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_130(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_63.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_131(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_64.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_132(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_65.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_133(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_66.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_134(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_67.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_135(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_68.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_136(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_69.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_137(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_70.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_138(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_71.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_139(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_72.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_140(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_73.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_141(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_74.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_142(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_75.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_143(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_76.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_144(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_77.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_145(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_78.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_146(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_79.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_147(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_80.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_148(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_81.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_149(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_82.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_150(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_83.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_151(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_84.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_152(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_85.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_153(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_86.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_154(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_87.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_155(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_88.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_156(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_89.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_157(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_90.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_158(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_91.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_159(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_92.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_160(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_93.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_161(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_94.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_162(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_95.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_163(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_96.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_164(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_97.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_165(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_98.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_166(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_99.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_167(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_100.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_168(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_101.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_169(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_102.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_170(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_103.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_171(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_104.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_172(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_105.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_173(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_106.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_174(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_107.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_175(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_108.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_176(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_109.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_177(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_110.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_178(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_111.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_179(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_112.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_180(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_113.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_181(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_114.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_182(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_115.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_183(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_116.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_184(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_117.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_185(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_118.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_186(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_119.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_187(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_120.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_188(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_121.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_189(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_122.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_190(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_123.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_191(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_124.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_192(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_125.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_193(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_126.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_194(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_127.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module MultiHotPriortyReductionTree(
  input  [5:0] io_dataInput_0, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_1, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_2, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_3, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_4, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_5, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_6, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_7, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_8, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_9, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_10, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_11, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_12, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_13, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_14, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_15, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_16, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_17, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_18, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_19, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_20, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_21, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_22, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_23, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_24, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_25, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_26, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_27, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_28, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_29, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_30, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_31, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_32, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_33, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_34, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_35, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_36, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_37, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_38, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_39, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_40, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_41, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_42, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_43, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_44, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_45, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_46, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_47, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_48, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_49, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_50, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_51, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_52, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_53, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_54, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_55, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_56, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_57, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_58, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_59, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_60, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_61, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_62, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_63, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_64, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_65, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_66, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_67, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_68, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_69, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_70, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_71, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_72, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_73, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_74, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_75, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_76, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_77, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_78, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_79, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_80, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_81, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_82, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_83, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_84, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_85, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_86, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_87, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_88, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_89, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_90, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_91, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_92, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_93, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_94, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_95, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_96, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_97, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_98, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_99, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_100, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_101, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_102, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_103, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_104, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_105, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_106, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_107, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_108, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_109, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_110, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_111, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_112, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_113, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_114, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_115, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_116, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_117, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_118, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_119, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_120, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_121, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_122, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_123, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_124, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_125, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_126, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_127, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_0, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_1, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_2, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_3, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_4, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_5, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_6, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_7, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_8, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_9, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_10, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_11, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_12, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_13, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_14, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_15, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_16, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_17, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_18, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_19, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_20, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_21, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_22, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_23, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_24, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_25, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_26, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_27, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_28, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_29, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_30, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_31, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_32, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_33, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_34, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_35, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_36, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_37, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_38, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_39, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_40, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_41, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_42, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_43, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_44, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_45, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_46, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_47, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_48, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_49, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_50, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_51, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_52, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_53, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_54, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_55, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_56, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_57, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_58, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_59, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_60, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_61, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_62, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_63, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_64, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_65, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_66, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_67, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_68, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_69, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_70, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_71, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_72, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_73, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_74, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_75, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_76, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_77, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_78, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_79, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_80, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_81, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_82, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_83, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_84, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_85, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_86, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_87, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_88, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_89, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_90, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_91, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_92, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_93, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_94, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_95, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_96, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_97, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_98, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_99, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_100, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_101, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_102, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_103, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_104, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_105, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_106, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_107, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_108, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_109, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_110, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_111, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_112, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_113, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_114, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_115, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_116, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_117, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_118, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_119, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_120, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_121, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_122, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_123, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_124, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_125, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_126, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_127, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  output [5:0] io_dataOutput, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  output       io_selectOutput // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
);
  wire  selectNodeOutputs_63 = io_selectInput_0 | io_selectInput_1; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_64 = io_selectInput_2 | io_selectInput_3; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_31 = selectNodeOutputs_63 | selectNodeOutputs_64; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_65 = io_selectInput_4 | io_selectInput_5; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_66 = io_selectInput_6 | io_selectInput_7; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_32 = selectNodeOutputs_65 | selectNodeOutputs_66; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_15 = selectNodeOutputs_31 | selectNodeOutputs_32; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_67 = io_selectInput_8 | io_selectInput_9; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_68 = io_selectInput_10 | io_selectInput_11; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_33 = selectNodeOutputs_67 | selectNodeOutputs_68; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_69 = io_selectInput_12 | io_selectInput_13; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_70 = io_selectInput_14 | io_selectInput_15; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_34 = selectNodeOutputs_69 | selectNodeOutputs_70; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_16 = selectNodeOutputs_33 | selectNodeOutputs_34; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_7 = selectNodeOutputs_15 | selectNodeOutputs_16; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_71 = io_selectInput_16 | io_selectInput_17; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_72 = io_selectInput_18 | io_selectInput_19; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_35 = selectNodeOutputs_71 | selectNodeOutputs_72; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_73 = io_selectInput_20 | io_selectInput_21; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_74 = io_selectInput_22 | io_selectInput_23; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_36 = selectNodeOutputs_73 | selectNodeOutputs_74; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_17 = selectNodeOutputs_35 | selectNodeOutputs_36; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_75 = io_selectInput_24 | io_selectInput_25; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_76 = io_selectInput_26 | io_selectInput_27; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_37 = selectNodeOutputs_75 | selectNodeOutputs_76; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_77 = io_selectInput_28 | io_selectInput_29; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_78 = io_selectInput_30 | io_selectInput_31; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_38 = selectNodeOutputs_77 | selectNodeOutputs_78; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_18 = selectNodeOutputs_37 | selectNodeOutputs_38; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_8 = selectNodeOutputs_17 | selectNodeOutputs_18; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_3 = selectNodeOutputs_7 | selectNodeOutputs_8; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_79 = io_selectInput_32 | io_selectInput_33; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_80 = io_selectInput_34 | io_selectInput_35; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_39 = selectNodeOutputs_79 | selectNodeOutputs_80; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_81 = io_selectInput_36 | io_selectInput_37; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_82 = io_selectInput_38 | io_selectInput_39; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_40 = selectNodeOutputs_81 | selectNodeOutputs_82; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_19 = selectNodeOutputs_39 | selectNodeOutputs_40; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_83 = io_selectInput_40 | io_selectInput_41; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_84 = io_selectInput_42 | io_selectInput_43; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_41 = selectNodeOutputs_83 | selectNodeOutputs_84; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_85 = io_selectInput_44 | io_selectInput_45; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_86 = io_selectInput_46 | io_selectInput_47; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_42 = selectNodeOutputs_85 | selectNodeOutputs_86; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_20 = selectNodeOutputs_41 | selectNodeOutputs_42; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_9 = selectNodeOutputs_19 | selectNodeOutputs_20; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_87 = io_selectInput_48 | io_selectInput_49; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_88 = io_selectInput_50 | io_selectInput_51; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_43 = selectNodeOutputs_87 | selectNodeOutputs_88; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_89 = io_selectInput_52 | io_selectInput_53; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_90 = io_selectInput_54 | io_selectInput_55; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_44 = selectNodeOutputs_89 | selectNodeOutputs_90; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_21 = selectNodeOutputs_43 | selectNodeOutputs_44; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_91 = io_selectInput_56 | io_selectInput_57; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_92 = io_selectInput_58 | io_selectInput_59; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_45 = selectNodeOutputs_91 | selectNodeOutputs_92; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_93 = io_selectInput_60 | io_selectInput_61; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_94 = io_selectInput_62 | io_selectInput_63; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_46 = selectNodeOutputs_93 | selectNodeOutputs_94; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_22 = selectNodeOutputs_45 | selectNodeOutputs_46; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_10 = selectNodeOutputs_21 | selectNodeOutputs_22; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_4 = selectNodeOutputs_9 | selectNodeOutputs_10; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_1 = selectNodeOutputs_3 | selectNodeOutputs_4; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_63 = io_selectInput_0 ? io_dataInput_0 : io_dataInput_1; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_64 = io_selectInput_2 ? io_dataInput_2 : io_dataInput_3; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_31 = selectNodeOutputs_63 ? dataNodeOutputs_63 : dataNodeOutputs_64; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_65 = io_selectInput_4 ? io_dataInput_4 : io_dataInput_5; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_66 = io_selectInput_6 ? io_dataInput_6 : io_dataInput_7; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_32 = selectNodeOutputs_65 ? dataNodeOutputs_65 : dataNodeOutputs_66; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_15 = selectNodeOutputs_31 ? dataNodeOutputs_31 : dataNodeOutputs_32; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_67 = io_selectInput_8 ? io_dataInput_8 : io_dataInput_9; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_68 = io_selectInput_10 ? io_dataInput_10 : io_dataInput_11; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_33 = selectNodeOutputs_67 ? dataNodeOutputs_67 : dataNodeOutputs_68; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_69 = io_selectInput_12 ? io_dataInput_12 : io_dataInput_13; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_70 = io_selectInput_14 ? io_dataInput_14 : io_dataInput_15; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_34 = selectNodeOutputs_69 ? dataNodeOutputs_69 : dataNodeOutputs_70; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_16 = selectNodeOutputs_33 ? dataNodeOutputs_33 : dataNodeOutputs_34; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_7 = selectNodeOutputs_15 ? dataNodeOutputs_15 : dataNodeOutputs_16; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_71 = io_selectInput_16 ? io_dataInput_16 : io_dataInput_17; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_72 = io_selectInput_18 ? io_dataInput_18 : io_dataInput_19; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_35 = selectNodeOutputs_71 ? dataNodeOutputs_71 : dataNodeOutputs_72; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_73 = io_selectInput_20 ? io_dataInput_20 : io_dataInput_21; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_74 = io_selectInput_22 ? io_dataInput_22 : io_dataInput_23; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_36 = selectNodeOutputs_73 ? dataNodeOutputs_73 : dataNodeOutputs_74; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_17 = selectNodeOutputs_35 ? dataNodeOutputs_35 : dataNodeOutputs_36; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_75 = io_selectInput_24 ? io_dataInput_24 : io_dataInput_25; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_76 = io_selectInput_26 ? io_dataInput_26 : io_dataInput_27; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_37 = selectNodeOutputs_75 ? dataNodeOutputs_75 : dataNodeOutputs_76; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_77 = io_selectInput_28 ? io_dataInput_28 : io_dataInput_29; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_78 = io_selectInput_30 ? io_dataInput_30 : io_dataInput_31; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_38 = selectNodeOutputs_77 ? dataNodeOutputs_77 : dataNodeOutputs_78; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_18 = selectNodeOutputs_37 ? dataNodeOutputs_37 : dataNodeOutputs_38; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_8 = selectNodeOutputs_17 ? dataNodeOutputs_17 : dataNodeOutputs_18; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_3 = selectNodeOutputs_7 ? dataNodeOutputs_7 : dataNodeOutputs_8; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_79 = io_selectInput_32 ? io_dataInput_32 : io_dataInput_33; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_80 = io_selectInput_34 ? io_dataInput_34 : io_dataInput_35; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_39 = selectNodeOutputs_79 ? dataNodeOutputs_79 : dataNodeOutputs_80; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_81 = io_selectInput_36 ? io_dataInput_36 : io_dataInput_37; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_82 = io_selectInput_38 ? io_dataInput_38 : io_dataInput_39; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_40 = selectNodeOutputs_81 ? dataNodeOutputs_81 : dataNodeOutputs_82; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_19 = selectNodeOutputs_39 ? dataNodeOutputs_39 : dataNodeOutputs_40; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_83 = io_selectInput_40 ? io_dataInput_40 : io_dataInput_41; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_84 = io_selectInput_42 ? io_dataInput_42 : io_dataInput_43; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_41 = selectNodeOutputs_83 ? dataNodeOutputs_83 : dataNodeOutputs_84; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_85 = io_selectInput_44 ? io_dataInput_44 : io_dataInput_45; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_86 = io_selectInput_46 ? io_dataInput_46 : io_dataInput_47; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_42 = selectNodeOutputs_85 ? dataNodeOutputs_85 : dataNodeOutputs_86; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_20 = selectNodeOutputs_41 ? dataNodeOutputs_41 : dataNodeOutputs_42; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_9 = selectNodeOutputs_19 ? dataNodeOutputs_19 : dataNodeOutputs_20; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_87 = io_selectInput_48 ? io_dataInput_48 : io_dataInput_49; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_88 = io_selectInput_50 ? io_dataInput_50 : io_dataInput_51; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_43 = selectNodeOutputs_87 ? dataNodeOutputs_87 : dataNodeOutputs_88; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_89 = io_selectInput_52 ? io_dataInput_52 : io_dataInput_53; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_90 = io_selectInput_54 ? io_dataInput_54 : io_dataInput_55; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_44 = selectNodeOutputs_89 ? dataNodeOutputs_89 : dataNodeOutputs_90; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_21 = selectNodeOutputs_43 ? dataNodeOutputs_43 : dataNodeOutputs_44; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_91 = io_selectInput_56 ? io_dataInput_56 : io_dataInput_57; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_92 = io_selectInput_58 ? io_dataInput_58 : io_dataInput_59; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_45 = selectNodeOutputs_91 ? dataNodeOutputs_91 : dataNodeOutputs_92; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_93 = io_selectInput_60 ? io_dataInput_60 : io_dataInput_61; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_94 = io_selectInput_62 ? io_dataInput_62 : io_dataInput_63; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_46 = selectNodeOutputs_93 ? dataNodeOutputs_93 : dataNodeOutputs_94; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_22 = selectNodeOutputs_45 ? dataNodeOutputs_45 : dataNodeOutputs_46; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_10 = selectNodeOutputs_21 ? dataNodeOutputs_21 : dataNodeOutputs_22; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_4 = selectNodeOutputs_9 ? dataNodeOutputs_9 : dataNodeOutputs_10; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_1 = selectNodeOutputs_3 ? dataNodeOutputs_3 : dataNodeOutputs_4; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_95 = io_selectInput_64 | io_selectInput_65; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_96 = io_selectInput_66 | io_selectInput_67; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_47 = selectNodeOutputs_95 | selectNodeOutputs_96; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_97 = io_selectInput_68 | io_selectInput_69; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_98 = io_selectInput_70 | io_selectInput_71; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_48 = selectNodeOutputs_97 | selectNodeOutputs_98; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_23 = selectNodeOutputs_47 | selectNodeOutputs_48; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_99 = io_selectInput_72 | io_selectInput_73; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_100 = io_selectInput_74 | io_selectInput_75; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_49 = selectNodeOutputs_99 | selectNodeOutputs_100; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_101 = io_selectInput_76 | io_selectInput_77; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_102 = io_selectInput_78 | io_selectInput_79; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_50 = selectNodeOutputs_101 | selectNodeOutputs_102; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_24 = selectNodeOutputs_49 | selectNodeOutputs_50; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_11 = selectNodeOutputs_23 | selectNodeOutputs_24; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_103 = io_selectInput_80 | io_selectInput_81; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_104 = io_selectInput_82 | io_selectInput_83; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_51 = selectNodeOutputs_103 | selectNodeOutputs_104; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_105 = io_selectInput_84 | io_selectInput_85; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_106 = io_selectInput_86 | io_selectInput_87; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_52 = selectNodeOutputs_105 | selectNodeOutputs_106; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_25 = selectNodeOutputs_51 | selectNodeOutputs_52; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_107 = io_selectInput_88 | io_selectInput_89; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_108 = io_selectInput_90 | io_selectInput_91; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_53 = selectNodeOutputs_107 | selectNodeOutputs_108; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_109 = io_selectInput_92 | io_selectInput_93; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_110 = io_selectInput_94 | io_selectInput_95; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_54 = selectNodeOutputs_109 | selectNodeOutputs_110; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_26 = selectNodeOutputs_53 | selectNodeOutputs_54; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_12 = selectNodeOutputs_25 | selectNodeOutputs_26; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_5 = selectNodeOutputs_11 | selectNodeOutputs_12; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_95 = io_selectInput_64 ? io_dataInput_64 : io_dataInput_65; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_96 = io_selectInput_66 ? io_dataInput_66 : io_dataInput_67; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_47 = selectNodeOutputs_95 ? dataNodeOutputs_95 : dataNodeOutputs_96; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_97 = io_selectInput_68 ? io_dataInput_68 : io_dataInput_69; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_98 = io_selectInput_70 ? io_dataInput_70 : io_dataInput_71; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_48 = selectNodeOutputs_97 ? dataNodeOutputs_97 : dataNodeOutputs_98; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_23 = selectNodeOutputs_47 ? dataNodeOutputs_47 : dataNodeOutputs_48; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_99 = io_selectInput_72 ? io_dataInput_72 : io_dataInput_73; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_100 = io_selectInput_74 ? io_dataInput_74 : io_dataInput_75; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_49 = selectNodeOutputs_99 ? dataNodeOutputs_99 : dataNodeOutputs_100; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_101 = io_selectInput_76 ? io_dataInput_76 : io_dataInput_77; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_102 = io_selectInput_78 ? io_dataInput_78 : io_dataInput_79; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_50 = selectNodeOutputs_101 ? dataNodeOutputs_101 : dataNodeOutputs_102; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_24 = selectNodeOutputs_49 ? dataNodeOutputs_49 : dataNodeOutputs_50; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_11 = selectNodeOutputs_23 ? dataNodeOutputs_23 : dataNodeOutputs_24; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_103 = io_selectInput_80 ? io_dataInput_80 : io_dataInput_81; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_104 = io_selectInput_82 ? io_dataInput_82 : io_dataInput_83; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_51 = selectNodeOutputs_103 ? dataNodeOutputs_103 : dataNodeOutputs_104; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_105 = io_selectInput_84 ? io_dataInput_84 : io_dataInput_85; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_106 = io_selectInput_86 ? io_dataInput_86 : io_dataInput_87; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_52 = selectNodeOutputs_105 ? dataNodeOutputs_105 : dataNodeOutputs_106; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_25 = selectNodeOutputs_51 ? dataNodeOutputs_51 : dataNodeOutputs_52; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_107 = io_selectInput_88 ? io_dataInput_88 : io_dataInput_89; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_108 = io_selectInput_90 ? io_dataInput_90 : io_dataInput_91; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_53 = selectNodeOutputs_107 ? dataNodeOutputs_107 : dataNodeOutputs_108; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_109 = io_selectInput_92 ? io_dataInput_92 : io_dataInput_93; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_110 = io_selectInput_94 ? io_dataInput_94 : io_dataInput_95; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_54 = selectNodeOutputs_109 ? dataNodeOutputs_109 : dataNodeOutputs_110; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_26 = selectNodeOutputs_53 ? dataNodeOutputs_53 : dataNodeOutputs_54; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_12 = selectNodeOutputs_25 ? dataNodeOutputs_25 : dataNodeOutputs_26; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_5 = selectNodeOutputs_11 ? dataNodeOutputs_11 : dataNodeOutputs_12; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_111 = io_selectInput_96 | io_selectInput_97; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_112 = io_selectInput_98 | io_selectInput_99; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_55 = selectNodeOutputs_111 | selectNodeOutputs_112; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_113 = io_selectInput_100 | io_selectInput_101; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_114 = io_selectInput_102 | io_selectInput_103; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_56 = selectNodeOutputs_113 | selectNodeOutputs_114; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_27 = selectNodeOutputs_55 | selectNodeOutputs_56; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_115 = io_selectInput_104 | io_selectInput_105; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_116 = io_selectInput_106 | io_selectInput_107; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_57 = selectNodeOutputs_115 | selectNodeOutputs_116; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_117 = io_selectInput_108 | io_selectInput_109; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_118 = io_selectInput_110 | io_selectInput_111; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_58 = selectNodeOutputs_117 | selectNodeOutputs_118; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_28 = selectNodeOutputs_57 | selectNodeOutputs_58; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_13 = selectNodeOutputs_27 | selectNodeOutputs_28; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_111 = io_selectInput_96 ? io_dataInput_96 : io_dataInput_97; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_112 = io_selectInput_98 ? io_dataInput_98 : io_dataInput_99; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_55 = selectNodeOutputs_111 ? dataNodeOutputs_111 : dataNodeOutputs_112; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_113 = io_selectInput_100 ? io_dataInput_100 : io_dataInput_101; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_114 = io_selectInput_102 ? io_dataInput_102 : io_dataInput_103; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_56 = selectNodeOutputs_113 ? dataNodeOutputs_113 : dataNodeOutputs_114; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_27 = selectNodeOutputs_55 ? dataNodeOutputs_55 : dataNodeOutputs_56; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_115 = io_selectInput_104 ? io_dataInput_104 : io_dataInput_105; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_116 = io_selectInput_106 ? io_dataInput_106 : io_dataInput_107; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_57 = selectNodeOutputs_115 ? dataNodeOutputs_115 : dataNodeOutputs_116; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_117 = io_selectInput_108 ? io_dataInput_108 : io_dataInput_109; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_118 = io_selectInput_110 ? io_dataInput_110 : io_dataInput_111; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_58 = selectNodeOutputs_117 ? dataNodeOutputs_117 : dataNodeOutputs_118; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_28 = selectNodeOutputs_57 ? dataNodeOutputs_57 : dataNodeOutputs_58; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_13 = selectNodeOutputs_27 ? dataNodeOutputs_27 : dataNodeOutputs_28; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_119 = io_selectInput_112 | io_selectInput_113; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_120 = io_selectInput_114 | io_selectInput_115; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_59 = selectNodeOutputs_119 | selectNodeOutputs_120; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_121 = io_selectInput_116 | io_selectInput_117; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_122 = io_selectInput_118 | io_selectInput_119; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_60 = selectNodeOutputs_121 | selectNodeOutputs_122; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_29 = selectNodeOutputs_59 | selectNodeOutputs_60; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_119 = io_selectInput_112 ? io_dataInput_112 : io_dataInput_113; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_120 = io_selectInput_114 ? io_dataInput_114 : io_dataInput_115; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_59 = selectNodeOutputs_119 ? dataNodeOutputs_119 : dataNodeOutputs_120; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_121 = io_selectInput_116 ? io_dataInput_116 : io_dataInput_117; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_122 = io_selectInput_118 ? io_dataInput_118 : io_dataInput_119; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_60 = selectNodeOutputs_121 ? dataNodeOutputs_121 : dataNodeOutputs_122; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_29 = selectNodeOutputs_59 ? dataNodeOutputs_59 : dataNodeOutputs_60; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_123 = io_selectInput_120 | io_selectInput_121; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_124 = io_selectInput_122 | io_selectInput_123; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_61 = selectNodeOutputs_123 | selectNodeOutputs_124; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_123 = io_selectInput_120 ? io_dataInput_120 : io_dataInput_121; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_124 = io_selectInput_122 ? io_dataInput_122 : io_dataInput_123; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_61 = selectNodeOutputs_123 ? dataNodeOutputs_123 : dataNodeOutputs_124; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_125 = io_selectInput_124 | io_selectInput_125; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_125 = io_selectInput_124 ? io_dataInput_124 : io_dataInput_125; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_126 = io_selectInput_126 ? io_dataInput_126 : io_dataInput_127; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_62 = selectNodeOutputs_125 ? dataNodeOutputs_125 : dataNodeOutputs_126; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_30 = selectNodeOutputs_61 ? dataNodeOutputs_61 : dataNodeOutputs_62; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_14 = selectNodeOutputs_29 ? dataNodeOutputs_29 : dataNodeOutputs_30; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_6 = selectNodeOutputs_13 ? dataNodeOutputs_13 : dataNodeOutputs_14; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_2 = selectNodeOutputs_5 ? dataNodeOutputs_5 : dataNodeOutputs_6; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_126 = io_selectInput_126 | io_selectInput_127; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_62 = selectNodeOutputs_125 | selectNodeOutputs_126; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_30 = selectNodeOutputs_61 | selectNodeOutputs_62; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_14 = selectNodeOutputs_29 | selectNodeOutputs_30; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_6 = selectNodeOutputs_13 | selectNodeOutputs_14; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_2 = selectNodeOutputs_5 | selectNodeOutputs_6; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  assign io_dataOutput = selectNodeOutputs_1 ? dataNodeOutputs_1 : dataNodeOutputs_2; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  assign io_selectOutput = selectNodeOutputs_1 | selectNodeOutputs_2; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
endmodule
module GraphicEngineVGA(
  input         clock,
  input         reset,
  input  [10:0] io_spriteXPosition_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_46, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_47, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_48, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_49, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_50, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_51, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_52, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_53, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_54, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_55, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_56, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_57, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_61, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_62, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_63, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_46, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_47, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_48, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_49, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_50, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_51, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_52, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_53, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_54, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_55, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_56, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_57, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_61, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_62, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_63, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_4, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_5, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_6, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_15, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_46, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_47, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_48, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_49, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_50, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_51, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_52, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_53, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_54, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_55, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_56, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_57, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_61, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_62, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_63, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_64, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_65, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_66, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_67, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_68, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_69, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_70, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_71, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_72, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_73, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_74, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_75, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_76, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_77, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_78, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_79, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_80, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_81, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_82, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_83, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_84, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_85, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_86, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_87, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_88, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_89, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_90, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_91, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_92, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_93, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_94, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_95, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_96, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_97, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_98, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_99, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_viewBoxX, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [8:0]  io_viewBoxY, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_newFrame, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_frameUpdateDone, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_missingFrameError, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_viewBoxOutOfRangeError, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaRed, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaBlue, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaGreen, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_Hsync, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_Vsync // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
`endif // RANDOMIZE_REG_INIT
  wire  backTileMemories_0_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_0_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_1_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_1_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_2_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_2_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_3_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_3_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_4_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_4_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_5_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_5_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_6_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_6_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_7_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_7_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_8_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_8_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_9_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_9_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_10_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_10_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_11_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_11_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_12_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_12_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_13_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_13_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_14_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_14_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_15_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_15_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_16_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_16_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_17_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_17_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_18_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_18_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_19_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_19_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_20_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_20_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_21_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_21_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_22_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_22_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_23_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_23_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_24_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_24_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_25_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_25_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_26_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_26_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_27_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_27_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_28_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_28_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_29_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_29_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_30_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_30_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_31_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_31_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_32_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_32_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_32_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_33_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_33_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_33_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_34_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_34_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_34_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_35_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_35_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_35_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_36_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_36_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_36_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_37_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_37_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_37_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_38_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_38_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_38_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_39_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_39_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_39_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_40_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_40_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_40_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_41_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_41_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_41_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_42_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_42_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_42_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_43_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_43_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_43_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_44_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_44_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_44_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_45_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_45_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_45_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_46_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_46_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_46_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_47_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_47_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_47_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_48_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_48_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_48_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_49_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_49_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_49_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_50_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_50_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_50_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_51_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_51_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_51_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_52_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_52_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_52_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_53_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_53_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_53_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_54_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_54_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_54_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_55_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_55_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_55_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_56_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_56_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_56_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_57_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_57_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_57_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_58_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_58_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_58_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_59_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_59_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_59_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_60_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_60_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_60_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_61_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_61_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_61_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_62_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_62_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_62_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_63_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_63_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_63_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backBufferMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [10:0] backBufferMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [5:0] backBufferMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire  backBufferMemory_io_writeEnable; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [5:0] backBufferMemory_io_dataWrite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire  backBufferShadowMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [10:0] backBufferShadowMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [5:0] backBufferShadowMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire  backBufferShadowMemory_io_writeEnable; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [5:0] backBufferShadowMemory_io_dataWrite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire  backBufferRestoreMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire [10:0] backBufferRestoreMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire [5:0] backBufferRestoreMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire  spriteMemories_0_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_0_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_1_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_1_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_2_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_2_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_3_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_3_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_4_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_4_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_5_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_5_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_6_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_6_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_7_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_7_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_8_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_8_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_9_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_9_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_10_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_10_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_11_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_11_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_12_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_12_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_13_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_13_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_14_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_14_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_15_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_15_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_16_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_16_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_17_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_17_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_18_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_18_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_19_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_19_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_20_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_20_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_21_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_21_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_22_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_22_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_23_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_23_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_24_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_24_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_25_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_25_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_26_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_26_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_27_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_27_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_28_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_28_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_29_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_29_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_30_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_30_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_31_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_31_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_32_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_32_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_32_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_33_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_33_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_33_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_34_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_34_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_34_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_35_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_35_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_35_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_36_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_36_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_36_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_37_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_37_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_37_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_38_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_38_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_38_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_39_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_39_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_39_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_40_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_40_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_40_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_41_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_41_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_41_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_42_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_42_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_42_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_43_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_43_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_43_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_44_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_44_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_44_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_45_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_45_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_45_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_46_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_46_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_46_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_47_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_47_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_47_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_48_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_48_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_48_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_49_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_49_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_49_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_50_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_50_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_50_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_51_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_51_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_51_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_52_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_52_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_52_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_53_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_53_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_53_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_54_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_54_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_54_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_55_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_55_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_55_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_56_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_56_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_56_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_57_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_57_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_57_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_58_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_58_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_58_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_59_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_59_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_59_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_60_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_60_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_60_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_61_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_61_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_61_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_62_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_62_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_62_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_63_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_63_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_63_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_64_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_64_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_64_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_65_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_65_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_65_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_66_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_66_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_66_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_67_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_67_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_67_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_68_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_68_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_68_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_69_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_69_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_69_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_70_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_70_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_70_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_71_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_71_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_71_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_72_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_72_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_72_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_73_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_73_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_73_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_74_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_74_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_74_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_75_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_75_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_75_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_76_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_76_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_76_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_77_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_77_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_77_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_78_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_78_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_78_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_79_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_79_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_79_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_80_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_80_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_80_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_81_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_81_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_81_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_82_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_82_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_82_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_83_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_83_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_83_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_84_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_84_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_84_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_85_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_85_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_85_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_86_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_86_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_86_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_87_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_87_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_87_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_88_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_88_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_88_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_89_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_89_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_89_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_90_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_90_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_90_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_91_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_91_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_91_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_92_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_92_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_92_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_93_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_93_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_93_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_94_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_94_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_94_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_95_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_95_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_95_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_96_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_96_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_96_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_97_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_97_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_97_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_98_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_98_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_98_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_99_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_99_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_99_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_100_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_100_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_100_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_101_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_101_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_101_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_102_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_102_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_102_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_103_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_103_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_103_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_104_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_104_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_104_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_105_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_105_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_105_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_106_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_106_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_106_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_107_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_107_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_107_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_108_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_108_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_108_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_109_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_109_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_109_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_110_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_110_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_110_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_111_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_111_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_111_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_112_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_112_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_112_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_113_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_113_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_113_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_114_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_114_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_114_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_115_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_115_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_115_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_116_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_116_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_116_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_117_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_117_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_117_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_118_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_118_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_118_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_119_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_119_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_119_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_120_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_120_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_120_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_121_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_121_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_121_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_122_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_122_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_122_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_123_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_123_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_123_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_124_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_124_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_124_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_125_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_125_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_125_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_126_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_126_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_126_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_127_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_127_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_127_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_64; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_65; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_66; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_67; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_68; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_69; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_70; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_71; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_72; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_73; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_74; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_75; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_76; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_77; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_78; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_79; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_80; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_81; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_82; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_83; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_84; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_85; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_86; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_87; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_88; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_89; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_90; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_91; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_92; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_93; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_94; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_95; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_96; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_97; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_98; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_99; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_100; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_101; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_102; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_103; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_104; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_105; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_106; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_107; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_108; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_109; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_110; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_111; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_112; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_113; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_114; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_115; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_116; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_117; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_118; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_119; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_120; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_121; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_122; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_123; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_124; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_125; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_126; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_127; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_64; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_65; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_66; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_67; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_68; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_69; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_70; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_71; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_72; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_73; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_74; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_75; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_76; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_77; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_78; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_79; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_80; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_81; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_82; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_83; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_84; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_85; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_86; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_87; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_88; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_89; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_90; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_91; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_92; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_93; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_94; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_95; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_96; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_97; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_98; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_99; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_100; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_101; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_102; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_103; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_104; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_105; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_106; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_107; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_108; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_109; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_110; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_111; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_112; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_113; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_114; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_115; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_116; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_117; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_118; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_119; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_120; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_121; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_122; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_123; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_124; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_125; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_126; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_127; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  reg [1:0] ScaleCounterReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
  reg [9:0] CounterXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
  reg [9:0] CounterYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
  wire  _T_2 = CounterYReg == 10'h20c; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 78:26]
  wire [9:0] _CounterYReg_T_1 = CounterYReg + 10'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 82:38]
  wire [9:0] _GEN_0 = CounterYReg == 10'h20c ? 10'h0 : _CounterYReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 78:131 79:23 82:23]
  wire [9:0] _CounterXReg_T_1 = CounterXReg + 10'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 85:36]
  wire  _GEN_4 = CounterXReg == 10'h31f & _T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129 71:15]
  wire [1:0] _ScaleCounterReg_T_1 = ScaleCounterReg + 2'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 88:42]
  wire  _GEN_8 = ScaleCounterReg == 2'h3 & _GEN_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 71:15 74:52]
  reg [11:0] backMemoryRestoreCounter; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
  wire  restoreEnabled = backMemoryRestoreCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:33]
  wire  run = restoreEnabled ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:70 209:9 213:9]
  wire  Hsync = CounterXReg >= 10'h290 & CounterXReg < 10'h2f0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 92:79]
  wire  Vsync = CounterYReg >= 10'h1ea & CounterYReg < 10'h1ec; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 93:79]
  reg  io_Hsync_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg [20:0] frameClockCount; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
  wire [20:0] _frameClockCount_T_2 = frameClockCount + 21'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 105:92]
  wire  preDisplayArea = frameClockCount >= 21'h199a1b; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 106:40]
  reg [10:0] spriteXPositionReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [9:0] spriteYPositionReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg  spriteVisibleReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_64; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_65; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_66; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_67; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_68; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_69; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_70; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_71; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_72; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_73; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_74; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_75; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_76; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_77; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_78; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_79; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_80; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_81; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_82; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_83; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_84; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_85; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_86; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_87; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_88; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_89; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_90; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_91; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_92; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_93; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_94; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_95; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_96; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_97; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_98; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_99; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_100; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_101; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_102; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_103; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_104; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_105; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_106; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_107; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_108; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_109; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_110; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_111; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_112; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_113; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_114; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_115; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_116; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_117; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_118; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_119; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_120; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_121; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_122; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_123; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_124; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_125; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_126; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_127; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  wire  _GEN_269 = io_newFrame ? 1'h0 : spriteVisibleReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_270 = io_newFrame ? 1'h0 : spriteVisibleReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_271 = io_newFrame ? 1'h0 : spriteVisibleReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_272 = io_newFrame ? io_spriteVisible_3 : spriteVisibleReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_273 = io_newFrame ? io_spriteVisible_4 : spriteVisibleReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_274 = io_newFrame ? io_spriteVisible_5 : spriteVisibleReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_275 = io_newFrame ? io_spriteVisible_6 : spriteVisibleReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_276 = io_newFrame ? io_spriteVisible_7 : spriteVisibleReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_277 = io_newFrame ? io_spriteVisible_8 : spriteVisibleReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_278 = io_newFrame ? io_spriteVisible_9 : spriteVisibleReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_279 = io_newFrame ? io_spriteVisible_10 : spriteVisibleReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_280 = io_newFrame ? io_spriteVisible_11 : spriteVisibleReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_281 = io_newFrame ? io_spriteVisible_12 : spriteVisibleReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_282 = io_newFrame ? io_spriteVisible_13 : spriteVisibleReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_283 = io_newFrame ? io_spriteVisible_14 : spriteVisibleReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_284 = io_newFrame ? io_spriteVisible_15 : spriteVisibleReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_285 = io_newFrame ? io_spriteVisible_16 : spriteVisibleReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_286 = io_newFrame ? io_spriteVisible_17 : spriteVisibleReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_287 = io_newFrame ? io_spriteVisible_18 : spriteVisibleReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_288 = io_newFrame ? io_spriteVisible_19 : spriteVisibleReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_289 = io_newFrame ? io_spriteVisible_20 : spriteVisibleReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_290 = io_newFrame ? io_spriteVisible_21 : spriteVisibleReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_291 = io_newFrame ? io_spriteVisible_22 : spriteVisibleReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_292 = io_newFrame ? io_spriteVisible_23 : spriteVisibleReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_293 = io_newFrame ? io_spriteVisible_24 : spriteVisibleReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_294 = io_newFrame ? io_spriteVisible_25 : spriteVisibleReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_295 = io_newFrame ? io_spriteVisible_26 : spriteVisibleReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_296 = io_newFrame ? io_spriteVisible_27 : spriteVisibleReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_297 = io_newFrame ? io_spriteVisible_28 : spriteVisibleReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_298 = io_newFrame ? io_spriteVisible_29 : spriteVisibleReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_299 = io_newFrame ? io_spriteVisible_30 : spriteVisibleReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_300 = io_newFrame ? io_spriteVisible_31 : spriteVisibleReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_301 = io_newFrame ? io_spriteVisible_32 : spriteVisibleReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_302 = io_newFrame ? io_spriteVisible_33 : spriteVisibleReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_303 = io_newFrame ? io_spriteVisible_34 : spriteVisibleReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_304 = io_newFrame ? io_spriteVisible_35 : spriteVisibleReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_305 = io_newFrame ? io_spriteVisible_36 : spriteVisibleReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_306 = io_newFrame ? io_spriteVisible_37 : spriteVisibleReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_307 = io_newFrame ? io_spriteVisible_38 : spriteVisibleReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_308 = io_newFrame ? io_spriteVisible_39 : spriteVisibleReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_309 = io_newFrame ? io_spriteVisible_40 : spriteVisibleReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_310 = io_newFrame ? io_spriteVisible_41 : spriteVisibleReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_311 = io_newFrame ? io_spriteVisible_42 : spriteVisibleReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_312 = io_newFrame ? io_spriteVisible_43 : spriteVisibleReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_313 = io_newFrame ? io_spriteVisible_44 : spriteVisibleReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_314 = io_newFrame ? io_spriteVisible_45 : spriteVisibleReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_315 = io_newFrame ? io_spriteVisible_46 : spriteVisibleReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_316 = io_newFrame ? io_spriteVisible_47 : spriteVisibleReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_317 = io_newFrame ? io_spriteVisible_48 : spriteVisibleReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_318 = io_newFrame ? io_spriteVisible_49 : spriteVisibleReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_319 = io_newFrame ? io_spriteVisible_50 : spriteVisibleReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_320 = io_newFrame ? io_spriteVisible_51 : spriteVisibleReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_321 = io_newFrame ? io_spriteVisible_52 : spriteVisibleReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_322 = io_newFrame ? io_spriteVisible_53 : spriteVisibleReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_323 = io_newFrame ? io_spriteVisible_54 : spriteVisibleReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_324 = io_newFrame ? io_spriteVisible_55 : spriteVisibleReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_325 = io_newFrame ? io_spriteVisible_56 : spriteVisibleReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_326 = io_newFrame ? io_spriteVisible_57 : spriteVisibleReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_327 = io_newFrame ? io_spriteVisible_58 : spriteVisibleReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_328 = io_newFrame ? io_spriteVisible_59 : spriteVisibleReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_329 = io_newFrame ? io_spriteVisible_60 : spriteVisibleReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_330 = io_newFrame ? io_spriteVisible_61 : spriteVisibleReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_331 = io_newFrame ? io_spriteVisible_62 : spriteVisibleReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_332 = io_newFrame ? io_spriteVisible_63 : spriteVisibleReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_333 = io_newFrame ? io_spriteVisible_64 : spriteVisibleReg_64; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_334 = io_newFrame ? io_spriteVisible_65 : spriteVisibleReg_65; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_335 = io_newFrame ? io_spriteVisible_66 : spriteVisibleReg_66; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_336 = io_newFrame ? io_spriteVisible_67 : spriteVisibleReg_67; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_337 = io_newFrame ? io_spriteVisible_68 : spriteVisibleReg_68; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_338 = io_newFrame ? io_spriteVisible_69 : spriteVisibleReg_69; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_339 = io_newFrame ? io_spriteVisible_70 : spriteVisibleReg_70; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_340 = io_newFrame ? io_spriteVisible_71 : spriteVisibleReg_71; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_341 = io_newFrame ? io_spriteVisible_72 : spriteVisibleReg_72; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_342 = io_newFrame ? io_spriteVisible_73 : spriteVisibleReg_73; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_343 = io_newFrame ? io_spriteVisible_74 : spriteVisibleReg_74; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_344 = io_newFrame ? io_spriteVisible_75 : spriteVisibleReg_75; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_345 = io_newFrame ? io_spriteVisible_76 : spriteVisibleReg_76; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_346 = io_newFrame ? io_spriteVisible_77 : spriteVisibleReg_77; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_347 = io_newFrame ? io_spriteVisible_78 : spriteVisibleReg_78; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_348 = io_newFrame ? io_spriteVisible_79 : spriteVisibleReg_79; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_349 = io_newFrame ? io_spriteVisible_80 : spriteVisibleReg_80; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_350 = io_newFrame ? io_spriteVisible_81 : spriteVisibleReg_81; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_351 = io_newFrame ? io_spriteVisible_82 : spriteVisibleReg_82; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_352 = io_newFrame ? io_spriteVisible_83 : spriteVisibleReg_83; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_353 = io_newFrame ? io_spriteVisible_84 : spriteVisibleReg_84; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_354 = io_newFrame ? io_spriteVisible_85 : spriteVisibleReg_85; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_355 = io_newFrame ? io_spriteVisible_86 : spriteVisibleReg_86; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_356 = io_newFrame ? io_spriteVisible_87 : spriteVisibleReg_87; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_357 = io_newFrame ? io_spriteVisible_88 : spriteVisibleReg_88; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_358 = io_newFrame ? io_spriteVisible_89 : spriteVisibleReg_89; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_359 = io_newFrame ? io_spriteVisible_90 : spriteVisibleReg_90; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_360 = io_newFrame ? io_spriteVisible_91 : spriteVisibleReg_91; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_361 = io_newFrame ? io_spriteVisible_92 : spriteVisibleReg_92; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_362 = io_newFrame ? io_spriteVisible_93 : spriteVisibleReg_93; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_363 = io_newFrame ? io_spriteVisible_94 : spriteVisibleReg_94; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_364 = io_newFrame ? io_spriteVisible_95 : spriteVisibleReg_95; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_365 = io_newFrame ? io_spriteVisible_96 : spriteVisibleReg_96; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_366 = io_newFrame ? io_spriteVisible_97 : spriteVisibleReg_97; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_367 = io_newFrame ? io_spriteVisible_98 : spriteVisibleReg_98; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_368 = io_newFrame ? io_spriteVisible_99 : spriteVisibleReg_99; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_369 = io_newFrame ? 1'h0 : spriteVisibleReg_100; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_370 = io_newFrame ? 1'h0 : spriteVisibleReg_101; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_371 = io_newFrame ? 1'h0 : spriteVisibleReg_102; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_372 = io_newFrame ? 1'h0 : spriteVisibleReg_103; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_373 = io_newFrame ? 1'h0 : spriteVisibleReg_104; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_374 = io_newFrame ? 1'h0 : spriteVisibleReg_105; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_375 = io_newFrame ? 1'h0 : spriteVisibleReg_106; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_376 = io_newFrame ? 1'h0 : spriteVisibleReg_107; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_377 = io_newFrame ? 1'h0 : spriteVisibleReg_108; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_378 = io_newFrame ? 1'h0 : spriteVisibleReg_109; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_379 = io_newFrame ? 1'h0 : spriteVisibleReg_110; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_380 = io_newFrame ? 1'h0 : spriteVisibleReg_111; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_381 = io_newFrame ? 1'h0 : spriteVisibleReg_112; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_382 = io_newFrame ? 1'h0 : spriteVisibleReg_113; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_383 = io_newFrame ? 1'h0 : spriteVisibleReg_114; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_384 = io_newFrame ? 1'h0 : spriteVisibleReg_115; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_385 = io_newFrame ? 1'h0 : spriteVisibleReg_116; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_386 = io_newFrame ? 1'h0 : spriteVisibleReg_117; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_387 = io_newFrame ? 1'h0 : spriteVisibleReg_118; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_388 = io_newFrame ? 1'h0 : spriteVisibleReg_119; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_389 = io_newFrame ? 1'h0 : spriteVisibleReg_120; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_390 = io_newFrame ? 1'h0 : spriteVisibleReg_121; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_391 = io_newFrame ? 1'h0 : spriteVisibleReg_122; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_392 = io_newFrame ? 1'h0 : spriteVisibleReg_123; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_393 = io_newFrame ? 1'h0 : spriteVisibleReg_124; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_394 = io_newFrame ? 1'h0 : spriteVisibleReg_125; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_395 = io_newFrame ? 1'h0 : spriteVisibleReg_126; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_396 = io_newFrame ? 1'h0 : spriteVisibleReg_127; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  reg  spriteScaleUpHorizontalReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpVerticalReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg [9:0] viewBoxXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
  reg [8:0] viewBoxYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
  reg  missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
  reg  viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
  wire [9:0] viewBoxXClipped = viewBoxXReg >= 10'h280 ? 10'h280 : viewBoxXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 137:28]
  wire [8:0] viewBoxYClipped = viewBoxYReg >= 9'h1e0 ? 9'h1e0 : viewBoxYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 138:28]
  wire [10:0] pixelXBack = CounterXReg + viewBoxXClipped; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 139:27]
  wire [9:0] _GEN_3292 = {{1'd0}, viewBoxYClipped}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 140:27]
  wire [10:0] pixelYBack = CounterYReg + _GEN_3292; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 140:27]
  wire  _GEN_1167 = viewBoxXReg > 10'h280 | viewBoxYReg > 9'h1e0 | viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 141:51 142:31 130:42]
  reg  newFrameStikyReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
  wire  _GEN_1168 = io_newFrame | newFrameStikyReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 148:21 149:22 147:33]
  reg  REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:16]
  wire  _GEN_1170 = newFrameStikyReg & io_newFrame | missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 154:41 155:26 128:37]
  wire [10:0] _backTileMemories_0_io_address_T_2 = 6'h20 * pixelYBack[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:75]
  wire [10:0] _GEN_3293 = {{6'd0}, pixelXBack[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:62]
  wire [11:0] _backTileMemories_0_io_address_T_3 = _GEN_3293 + _backTileMemories_0_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:62]
  reg [6:0] backTileMemoryDataRead_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [11:0] backMemoryCopyCounter; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
  wire  _T_7 = backMemoryCopyCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 187:32]
  wire [11:0] _backMemoryCopyCounter_T_1 = backMemoryCopyCounter + 12'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 188:54]
  wire  copyEnabled = preDisplayArea & _T_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23 198:17]
  reg  copyEnabledReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 200:31]
  wire [11:0] _backMemoryRestoreCounter_T_1 = backMemoryRestoreCounter + 12'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 206:58]
  reg [10:0] backBufferShadowMemory_io_address_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:67]
  wire [10:0] _backBufferShadowMemory_io_address_T_2 = copyEnabled ? backMemoryCopyCounter[10:0] : 11'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:105]
  reg  backBufferShadowMemory_io_writeEnable_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:71]
  reg [10:0] backBufferMemory_io_address_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:61]
  wire [11:0] _backBufferMemory_io_address_T_3 = 6'h28 * pixelYBack[10:5]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:130]
  wire [11:0] _GEN_3357 = {{6'd0}, pixelXBack[10:5]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:117]
  wire [12:0] _backBufferMemory_io_address_T_4 = _GEN_3357 + _backBufferMemory_io_address_T_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:117]
  wire [12:0] _backBufferMemory_io_address_T_5 = copyEnabledReg ? {{2'd0}, backBufferMemory_io_address_REG} :
    _backBufferMemory_io_address_T_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:37]
  reg [5:0] fullBackgroundColor_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:56]
  wire [6:0] _GEN_1181 = 6'h1 == fullBackgroundColor_REG ? backTileMemoryDataRead_1_REG : backTileMemoryDataRead_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1182 = 6'h2 == fullBackgroundColor_REG ? backTileMemoryDataRead_2_REG : _GEN_1181; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1183 = 6'h3 == fullBackgroundColor_REG ? backTileMemoryDataRead_3_REG : _GEN_1182; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1184 = 6'h4 == fullBackgroundColor_REG ? backTileMemoryDataRead_4_REG : _GEN_1183; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1185 = 6'h5 == fullBackgroundColor_REG ? backTileMemoryDataRead_5_REG : _GEN_1184; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1186 = 6'h6 == fullBackgroundColor_REG ? backTileMemoryDataRead_6_REG : _GEN_1185; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1187 = 6'h7 == fullBackgroundColor_REG ? backTileMemoryDataRead_7_REG : _GEN_1186; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1188 = 6'h8 == fullBackgroundColor_REG ? backTileMemoryDataRead_8_REG : _GEN_1187; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1189 = 6'h9 == fullBackgroundColor_REG ? backTileMemoryDataRead_9_REG : _GEN_1188; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1190 = 6'ha == fullBackgroundColor_REG ? backTileMemoryDataRead_10_REG : _GEN_1189; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1191 = 6'hb == fullBackgroundColor_REG ? backTileMemoryDataRead_11_REG : _GEN_1190; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1192 = 6'hc == fullBackgroundColor_REG ? backTileMemoryDataRead_12_REG : _GEN_1191; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1193 = 6'hd == fullBackgroundColor_REG ? backTileMemoryDataRead_13_REG : _GEN_1192; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1194 = 6'he == fullBackgroundColor_REG ? backTileMemoryDataRead_14_REG : _GEN_1193; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1195 = 6'hf == fullBackgroundColor_REG ? backTileMemoryDataRead_15_REG : _GEN_1194; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1196 = 6'h10 == fullBackgroundColor_REG ? backTileMemoryDataRead_16_REG : _GEN_1195; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1197 = 6'h11 == fullBackgroundColor_REG ? backTileMemoryDataRead_17_REG : _GEN_1196; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1198 = 6'h12 == fullBackgroundColor_REG ? backTileMemoryDataRead_18_REG : _GEN_1197; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1199 = 6'h13 == fullBackgroundColor_REG ? backTileMemoryDataRead_19_REG : _GEN_1198; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1200 = 6'h14 == fullBackgroundColor_REG ? backTileMemoryDataRead_20_REG : _GEN_1199; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1201 = 6'h15 == fullBackgroundColor_REG ? backTileMemoryDataRead_21_REG : _GEN_1200; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1202 = 6'h16 == fullBackgroundColor_REG ? backTileMemoryDataRead_22_REG : _GEN_1201; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1203 = 6'h17 == fullBackgroundColor_REG ? backTileMemoryDataRead_23_REG : _GEN_1202; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1204 = 6'h18 == fullBackgroundColor_REG ? backTileMemoryDataRead_24_REG : _GEN_1203; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1205 = 6'h19 == fullBackgroundColor_REG ? backTileMemoryDataRead_25_REG : _GEN_1204; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1206 = 6'h1a == fullBackgroundColor_REG ? backTileMemoryDataRead_26_REG : _GEN_1205; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1207 = 6'h1b == fullBackgroundColor_REG ? backTileMemoryDataRead_27_REG : _GEN_1206; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1208 = 6'h1c == fullBackgroundColor_REG ? backTileMemoryDataRead_28_REG : _GEN_1207; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1209 = 6'h1d == fullBackgroundColor_REG ? backTileMemoryDataRead_29_REG : _GEN_1208; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1210 = 6'h1e == fullBackgroundColor_REG ? backTileMemoryDataRead_30_REG : _GEN_1209; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1211 = 6'h1f == fullBackgroundColor_REG ? backTileMemoryDataRead_31_REG : _GEN_1210; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1212 = 6'h20 == fullBackgroundColor_REG ? backTileMemoryDataRead_32_REG : _GEN_1211; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1213 = 6'h21 == fullBackgroundColor_REG ? backTileMemoryDataRead_33_REG : _GEN_1212; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1214 = 6'h22 == fullBackgroundColor_REG ? backTileMemoryDataRead_34_REG : _GEN_1213; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1215 = 6'h23 == fullBackgroundColor_REG ? backTileMemoryDataRead_35_REG : _GEN_1214; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1216 = 6'h24 == fullBackgroundColor_REG ? backTileMemoryDataRead_36_REG : _GEN_1215; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1217 = 6'h25 == fullBackgroundColor_REG ? backTileMemoryDataRead_37_REG : _GEN_1216; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1218 = 6'h26 == fullBackgroundColor_REG ? backTileMemoryDataRead_38_REG : _GEN_1217; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1219 = 6'h27 == fullBackgroundColor_REG ? backTileMemoryDataRead_39_REG : _GEN_1218; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1220 = 6'h28 == fullBackgroundColor_REG ? backTileMemoryDataRead_40_REG : _GEN_1219; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1221 = 6'h29 == fullBackgroundColor_REG ? backTileMemoryDataRead_41_REG : _GEN_1220; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1222 = 6'h2a == fullBackgroundColor_REG ? backTileMemoryDataRead_42_REG : _GEN_1221; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1223 = 6'h2b == fullBackgroundColor_REG ? backTileMemoryDataRead_43_REG : _GEN_1222; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1224 = 6'h2c == fullBackgroundColor_REG ? backTileMemoryDataRead_44_REG : _GEN_1223; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1225 = 6'h2d == fullBackgroundColor_REG ? backTileMemoryDataRead_45_REG : _GEN_1224; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1226 = 6'h2e == fullBackgroundColor_REG ? backTileMemoryDataRead_46_REG : _GEN_1225; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1227 = 6'h2f == fullBackgroundColor_REG ? backTileMemoryDataRead_47_REG : _GEN_1226; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1228 = 6'h30 == fullBackgroundColor_REG ? backTileMemoryDataRead_48_REG : _GEN_1227; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1229 = 6'h31 == fullBackgroundColor_REG ? backTileMemoryDataRead_49_REG : _GEN_1228; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1230 = 6'h32 == fullBackgroundColor_REG ? backTileMemoryDataRead_50_REG : _GEN_1229; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1231 = 6'h33 == fullBackgroundColor_REG ? backTileMemoryDataRead_51_REG : _GEN_1230; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1232 = 6'h34 == fullBackgroundColor_REG ? backTileMemoryDataRead_52_REG : _GEN_1231; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1233 = 6'h35 == fullBackgroundColor_REG ? backTileMemoryDataRead_53_REG : _GEN_1232; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1234 = 6'h36 == fullBackgroundColor_REG ? backTileMemoryDataRead_54_REG : _GEN_1233; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1235 = 6'h37 == fullBackgroundColor_REG ? backTileMemoryDataRead_55_REG : _GEN_1234; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1236 = 6'h38 == fullBackgroundColor_REG ? backTileMemoryDataRead_56_REG : _GEN_1235; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1237 = 6'h39 == fullBackgroundColor_REG ? backTileMemoryDataRead_57_REG : _GEN_1236; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1238 = 6'h3a == fullBackgroundColor_REG ? backTileMemoryDataRead_58_REG : _GEN_1237; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1239 = 6'h3b == fullBackgroundColor_REG ? backTileMemoryDataRead_59_REG : _GEN_1238; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1240 = 6'h3c == fullBackgroundColor_REG ? backTileMemoryDataRead_60_REG : _GEN_1239; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1241 = 6'h3d == fullBackgroundColor_REG ? backTileMemoryDataRead_61_REG : _GEN_1240; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_1242 = 6'h3e == fullBackgroundColor_REG ? backTileMemoryDataRead_62_REG : _GEN_1241; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] fullBackgroundColor = 6'h3f == fullBackgroundColor_REG ? backTileMemoryDataRead_63_REG : _GEN_1242; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  reg [5:0] pixelColorBack; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 245:31]
  wire [10:0] _inSpriteXValue_T_1 = {1'h0,CounterXReg}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:47]
  wire [11:0] inSpriteXValue = $signed(_inSpriteXValue_T_1) - 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_0 = $signed(inSpriteXValue) >= 12'sh0 & $signed(inSpriteXValue) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1250 = {{1{inSpriteXValue[11]}},inSpriteXValue}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _inSpriteYValue_T_1 = {1'h0,CounterYReg}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:47]
  wire [11:0] inSpriteYValue = $signed(_inSpriteYValue_T_1) - 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_0 = inSpriteYValue[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_0 = $signed(inSpriteYPreScaled_0) >= 11'sh0 & $signed(inSpriteYPreScaled_0) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1258 = {{1{inSpriteYPreScaled_0[10]}},inSpriteYPreScaled_0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_3 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_3); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_3 = $signed(inSpriteXValue_3) >= 12'sh0 & $signed(inSpriteXValue_3) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1298 = {{1{inSpriteXValue_3[11]}},inSpriteXValue_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3361 = {{1{spriteYPositionReg_3[9]}},spriteYPositionReg_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_3 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3361); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_3 = inSpriteYValue_3[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_3 = $signed(inSpriteYPreScaled_3) >= 11'sh0 & $signed(inSpriteYPreScaled_3) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1306 = {{1{inSpriteYPreScaled_3[10]}},inSpriteYPreScaled_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_7 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_7); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_7 = $signed(inSpriteXValue_7) >= 12'sh0 & $signed(inSpriteXValue_7) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1362 = {{1{inSpriteXValue_7[11]}},inSpriteXValue_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3366 = {{1{spriteYPositionReg_7[9]}},spriteYPositionReg_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_7 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3366); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_7 = inSpriteYValue_7[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_7 = $signed(inSpriteYPreScaled_7) >= 11'sh0 & $signed(inSpriteYPreScaled_7) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1370 = {{1{inSpriteYPreScaled_7[10]}},inSpriteYPreScaled_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_8 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_8); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_8 = $signed(inSpriteXValue_8) >= 12'sh0 & $signed(inSpriteXValue_8) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1378 = {{1{inSpriteXValue_8[11]}},inSpriteXValue_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3368 = {{1{spriteYPositionReg_8[9]}},spriteYPositionReg_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_8 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3368); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_8 = inSpriteYValue_8[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_8 = $signed(inSpriteYPreScaled_8) >= 11'sh0 & $signed(inSpriteYPreScaled_8) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1386 = {{1{inSpriteYPreScaled_8[10]}},inSpriteYPreScaled_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_9 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_9); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_9 = $signed(inSpriteXValue_9) >= 12'sh0 & $signed(inSpriteXValue_9) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1394 = {{1{inSpriteXValue_9[11]}},inSpriteXValue_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3370 = {{1{spriteYPositionReg_9[9]}},spriteYPositionReg_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_9 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3370); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_9 = inSpriteYValue_9[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_9 = $signed(inSpriteYPreScaled_9) >= 11'sh0 & $signed(inSpriteYPreScaled_9) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1402 = {{1{inSpriteYPreScaled_9[10]}},inSpriteYPreScaled_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_10 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_10); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_10 = $signed(inSpriteXValue_10) >= 12'sh0 & $signed(inSpriteXValue_10) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1410 = {{1{inSpriteXValue_10[11]}},inSpriteXValue_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3372 = {{1{spriteYPositionReg_10[9]}},spriteYPositionReg_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_10 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3372); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_10 = inSpriteYValue_10[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_10 = $signed(inSpriteYPreScaled_10) >= 11'sh0 & $signed(inSpriteYPreScaled_10) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1418 = {{1{inSpriteYPreScaled_10[10]}},inSpriteYPreScaled_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_11 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_11); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_11 = $signed(inSpriteXValue_11) >= 12'sh0 & $signed(inSpriteXValue_11) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1426 = {{1{inSpriteXValue_11[11]}},inSpriteXValue_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3374 = {{1{spriteYPositionReg_11[9]}},spriteYPositionReg_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_11 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3374); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_11 = inSpriteYValue_11[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_11 = $signed(inSpriteYPreScaled_11) >= 11'sh0 & $signed(inSpriteYPreScaled_11) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1434 = {{1{inSpriteYPreScaled_11[10]}},inSpriteYPreScaled_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_12 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_12); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_12 = $signed(inSpriteXValue_12) >= 12'sh0 & $signed(inSpriteXValue_12) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1442 = {{1{inSpriteXValue_12[11]}},inSpriteXValue_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3376 = {{1{spriteYPositionReg_12[9]}},spriteYPositionReg_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_12 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3376); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_12 = inSpriteYValue_12[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_12 = $signed(inSpriteYPreScaled_12) >= 11'sh0 & $signed(inSpriteYPreScaled_12) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1450 = {{1{inSpriteYPreScaled_12[10]}},inSpriteYPreScaled_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_13 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_13); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_13 = $signed(inSpriteXValue_13) >= 12'sh0 & $signed(inSpriteXValue_13) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1458 = {{1{inSpriteXValue_13[11]}},inSpriteXValue_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3378 = {{1{spriteYPositionReg_13[9]}},spriteYPositionReg_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_13 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3378); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_13 = inSpriteYValue_13[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_13 = $signed(inSpriteYPreScaled_13) >= 11'sh0 & $signed(inSpriteYPreScaled_13) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1466 = {{1{inSpriteYPreScaled_13[10]}},inSpriteYPreScaled_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_14 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_14); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_14 = $signed(inSpriteXValue_14) >= 12'sh0 & $signed(inSpriteXValue_14) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1474 = {{1{inSpriteXValue_14[11]}},inSpriteXValue_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3380 = {{1{spriteYPositionReg_14[9]}},spriteYPositionReg_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_14 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3380); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_14 = inSpriteYValue_14[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_14 = $signed(inSpriteYPreScaled_14) >= 11'sh0 & $signed(inSpriteYPreScaled_14) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1482 = {{1{inSpriteYPreScaled_14[10]}},inSpriteYPreScaled_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_16 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_16); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_16_T = $signed(inSpriteXValue_16) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_16_T_4 = inSpriteXValue_16[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_16_T_8 = _inSpriteHorizontal_16_T & $signed(inSpriteXValue_16) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_16_T_5 = {$signed(inSpriteXValue_16), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_16_T_14 = _inSpriteHorizontal_16_T & $signed(inSpriteXValue_16) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1504 = spriteScaleUpHorizontalReg_16 ? $signed({{2{_inSpriteX_16_T_4[10]}},_inSpriteX_16_T_4}) :
    $signed(_inSpriteX_16_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1505 = spriteScaleUpHorizontalReg_16 ? _inSpriteHorizontal_16_T_8 : _inSpriteHorizontal_16_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1506 = ~spriteScaleUpHorizontalReg_16 ? $signed({{1{inSpriteXValue_16[11]}},inSpriteXValue_16}) :
    $signed(_GEN_1504); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_16 = ~spriteScaleUpHorizontalReg_16 ? $signed(inSpriteXValue_16) >= 12'sh0 & $signed(
    inSpriteXValue_16) < 12'sh20 : _GEN_1505; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3383 = {{1{spriteYPositionReg_16[9]}},spriteYPositionReg_16}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_16 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3383); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_16 = inSpriteYValue_16[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_16_T = $signed(inSpriteYPreScaled_16) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_16_T_4 = inSpriteYPreScaled_16[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_16_T_8 = _inSpriteVertical_16_T & $signed(inSpriteYPreScaled_16) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_16_T_5 = {$signed(inSpriteYPreScaled_16), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_16_T_14 = _inSpriteVertical_16_T & $signed(inSpriteYPreScaled_16) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1512 = spriteScaleUpVerticalReg_16 ? $signed({{2{_inSpriteY_16_T_4[9]}},_inSpriteY_16_T_4}) :
    $signed(_inSpriteY_16_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1513 = spriteScaleUpVerticalReg_16 ? _inSpriteVertical_16_T_8 : _inSpriteVertical_16_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1514 = ~spriteScaleUpVerticalReg_16 ? $signed({{1{inSpriteYPreScaled_16[10]}},inSpriteYPreScaled_16})
     : $signed(_GEN_1512); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_16 = ~spriteScaleUpVerticalReg_16 ? $signed(inSpriteYPreScaled_16) >= 11'sh0 & $signed(
    inSpriteYPreScaled_16) < 11'sh20 : _GEN_1513; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_17 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_17); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_17_T = $signed(inSpriteXValue_17) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_17_T_4 = inSpriteXValue_17[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_17_T_8 = _inSpriteHorizontal_17_T & $signed(inSpriteXValue_17) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_17_T_5 = {$signed(inSpriteXValue_17), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_17_T_14 = _inSpriteHorizontal_17_T & $signed(inSpriteXValue_17) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1520 = spriteScaleUpHorizontalReg_17 ? $signed({{2{_inSpriteX_17_T_4[10]}},_inSpriteX_17_T_4}) :
    $signed(_inSpriteX_17_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1521 = spriteScaleUpHorizontalReg_17 ? _inSpriteHorizontal_17_T_8 : _inSpriteHorizontal_17_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1522 = ~spriteScaleUpHorizontalReg_17 ? $signed({{1{inSpriteXValue_17[11]}},inSpriteXValue_17}) :
    $signed(_GEN_1520); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_17 = ~spriteScaleUpHorizontalReg_17 ? $signed(inSpriteXValue_17) >= 12'sh0 & $signed(
    inSpriteXValue_17) < 12'sh20 : _GEN_1521; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3385 = {{1{spriteYPositionReg_17[9]}},spriteYPositionReg_17}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_17 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3385); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_17 = inSpriteYValue_17[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_17_T = $signed(inSpriteYPreScaled_17) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_17_T_4 = inSpriteYPreScaled_17[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_17_T_8 = _inSpriteVertical_17_T & $signed(inSpriteYPreScaled_17) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_17_T_5 = {$signed(inSpriteYPreScaled_17), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_17_T_14 = _inSpriteVertical_17_T & $signed(inSpriteYPreScaled_17) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1528 = spriteScaleUpVerticalReg_17 ? $signed({{2{_inSpriteY_17_T_4[9]}},_inSpriteY_17_T_4}) :
    $signed(_inSpriteY_17_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1529 = spriteScaleUpVerticalReg_17 ? _inSpriteVertical_17_T_8 : _inSpriteVertical_17_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1530 = ~spriteScaleUpVerticalReg_17 ? $signed({{1{inSpriteYPreScaled_17[10]}},inSpriteYPreScaled_17})
     : $signed(_GEN_1528); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_17 = ~spriteScaleUpVerticalReg_17 ? $signed(inSpriteYPreScaled_17) >= 11'sh0 & $signed(
    inSpriteYPreScaled_17) < 11'sh20 : _GEN_1529; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_18 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_18); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_18_T = $signed(inSpriteXValue_18) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_18_T_4 = inSpriteXValue_18[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_18_T_8 = _inSpriteHorizontal_18_T & $signed(inSpriteXValue_18) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_18_T_5 = {$signed(inSpriteXValue_18), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_18_T_14 = _inSpriteHorizontal_18_T & $signed(inSpriteXValue_18) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1536 = spriteScaleUpHorizontalReg_18 ? $signed({{2{_inSpriteX_18_T_4[10]}},_inSpriteX_18_T_4}) :
    $signed(_inSpriteX_18_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1537 = spriteScaleUpHorizontalReg_18 ? _inSpriteHorizontal_18_T_8 : _inSpriteHorizontal_18_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1538 = ~spriteScaleUpHorizontalReg_18 ? $signed({{1{inSpriteXValue_18[11]}},inSpriteXValue_18}) :
    $signed(_GEN_1536); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_18 = ~spriteScaleUpHorizontalReg_18 ? $signed(inSpriteXValue_18) >= 12'sh0 & $signed(
    inSpriteXValue_18) < 12'sh20 : _GEN_1537; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3387 = {{1{spriteYPositionReg_18[9]}},spriteYPositionReg_18}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_18 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3387); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_18 = inSpriteYValue_18[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_18_T = $signed(inSpriteYPreScaled_18) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_18_T_4 = inSpriteYPreScaled_18[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_18_T_8 = _inSpriteVertical_18_T & $signed(inSpriteYPreScaled_18) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_18_T_5 = {$signed(inSpriteYPreScaled_18), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_18_T_14 = _inSpriteVertical_18_T & $signed(inSpriteYPreScaled_18) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1544 = spriteScaleUpVerticalReg_18 ? $signed({{2{_inSpriteY_18_T_4[9]}},_inSpriteY_18_T_4}) :
    $signed(_inSpriteY_18_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1545 = spriteScaleUpVerticalReg_18 ? _inSpriteVertical_18_T_8 : _inSpriteVertical_18_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1546 = ~spriteScaleUpVerticalReg_18 ? $signed({{1{inSpriteYPreScaled_18[10]}},inSpriteYPreScaled_18})
     : $signed(_GEN_1544); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_18 = ~spriteScaleUpVerticalReg_18 ? $signed(inSpriteYPreScaled_18) >= 11'sh0 & $signed(
    inSpriteYPreScaled_18) < 11'sh20 : _GEN_1545; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_19 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_19); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_19_T = $signed(inSpriteXValue_19) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_19_T_4 = inSpriteXValue_19[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_19_T_8 = _inSpriteHorizontal_19_T & $signed(inSpriteXValue_19) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_19_T_5 = {$signed(inSpriteXValue_19), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_19_T_14 = _inSpriteHorizontal_19_T & $signed(inSpriteXValue_19) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1552 = spriteScaleUpHorizontalReg_19 ? $signed({{2{_inSpriteX_19_T_4[10]}},_inSpriteX_19_T_4}) :
    $signed(_inSpriteX_19_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1553 = spriteScaleUpHorizontalReg_19 ? _inSpriteHorizontal_19_T_8 : _inSpriteHorizontal_19_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1554 = ~spriteScaleUpHorizontalReg_19 ? $signed({{1{inSpriteXValue_19[11]}},inSpriteXValue_19}) :
    $signed(_GEN_1552); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_19 = ~spriteScaleUpHorizontalReg_19 ? $signed(inSpriteXValue_19) >= 12'sh0 & $signed(
    inSpriteXValue_19) < 12'sh20 : _GEN_1553; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3389 = {{1{spriteYPositionReg_19[9]}},spriteYPositionReg_19}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_19 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3389); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_19 = inSpriteYValue_19[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_19_T = $signed(inSpriteYPreScaled_19) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_19_T_4 = inSpriteYPreScaled_19[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_19_T_8 = _inSpriteVertical_19_T & $signed(inSpriteYPreScaled_19) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_19_T_5 = {$signed(inSpriteYPreScaled_19), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_19_T_14 = _inSpriteVertical_19_T & $signed(inSpriteYPreScaled_19) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1560 = spriteScaleUpVerticalReg_19 ? $signed({{2{_inSpriteY_19_T_4[9]}},_inSpriteY_19_T_4}) :
    $signed(_inSpriteY_19_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1561 = spriteScaleUpVerticalReg_19 ? _inSpriteVertical_19_T_8 : _inSpriteVertical_19_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1562 = ~spriteScaleUpVerticalReg_19 ? $signed({{1{inSpriteYPreScaled_19[10]}},inSpriteYPreScaled_19})
     : $signed(_GEN_1560); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_19 = ~spriteScaleUpVerticalReg_19 ? $signed(inSpriteYPreScaled_19) >= 11'sh0 & $signed(
    inSpriteYPreScaled_19) < 11'sh20 : _GEN_1561; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_20 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_20); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_20_T = $signed(inSpriteXValue_20) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_20_T_4 = inSpriteXValue_20[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_20_T_8 = _inSpriteHorizontal_20_T & $signed(inSpriteXValue_20) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_20_T_5 = {$signed(inSpriteXValue_20), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_20_T_14 = _inSpriteHorizontal_20_T & $signed(inSpriteXValue_20) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1568 = spriteScaleUpHorizontalReg_20 ? $signed({{2{_inSpriteX_20_T_4[10]}},_inSpriteX_20_T_4}) :
    $signed(_inSpriteX_20_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1569 = spriteScaleUpHorizontalReg_20 ? _inSpriteHorizontal_20_T_8 : _inSpriteHorizontal_20_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1570 = ~spriteScaleUpHorizontalReg_20 ? $signed({{1{inSpriteXValue_20[11]}},inSpriteXValue_20}) :
    $signed(_GEN_1568); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_20 = ~spriteScaleUpHorizontalReg_20 ? $signed(inSpriteXValue_20) >= 12'sh0 & $signed(
    inSpriteXValue_20) < 12'sh20 : _GEN_1569; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3391 = {{1{spriteYPositionReg_20[9]}},spriteYPositionReg_20}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_20 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3391); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_20 = inSpriteYValue_20[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_20_T = $signed(inSpriteYPreScaled_20) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_20_T_4 = inSpriteYPreScaled_20[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_20_T_8 = _inSpriteVertical_20_T & $signed(inSpriteYPreScaled_20) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_20_T_5 = {$signed(inSpriteYPreScaled_20), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_20_T_14 = _inSpriteVertical_20_T & $signed(inSpriteYPreScaled_20) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1576 = spriteScaleUpVerticalReg_20 ? $signed({{2{_inSpriteY_20_T_4[9]}},_inSpriteY_20_T_4}) :
    $signed(_inSpriteY_20_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1577 = spriteScaleUpVerticalReg_20 ? _inSpriteVertical_20_T_8 : _inSpriteVertical_20_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1578 = ~spriteScaleUpVerticalReg_20 ? $signed({{1{inSpriteYPreScaled_20[10]}},inSpriteYPreScaled_20})
     : $signed(_GEN_1576); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_20 = ~spriteScaleUpVerticalReg_20 ? $signed(inSpriteYPreScaled_20) >= 11'sh0 & $signed(
    inSpriteYPreScaled_20) < 11'sh20 : _GEN_1577; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_21 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_21); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_21_T = $signed(inSpriteXValue_21) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_21_T_4 = inSpriteXValue_21[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_21_T_8 = _inSpriteHorizontal_21_T & $signed(inSpriteXValue_21) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_21_T_5 = {$signed(inSpriteXValue_21), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_21_T_14 = _inSpriteHorizontal_21_T & $signed(inSpriteXValue_21) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1584 = spriteScaleUpHorizontalReg_21 ? $signed({{2{_inSpriteX_21_T_4[10]}},_inSpriteX_21_T_4}) :
    $signed(_inSpriteX_21_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1585 = spriteScaleUpHorizontalReg_21 ? _inSpriteHorizontal_21_T_8 : _inSpriteHorizontal_21_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1586 = ~spriteScaleUpHorizontalReg_21 ? $signed({{1{inSpriteXValue_21[11]}},inSpriteXValue_21}) :
    $signed(_GEN_1584); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_21 = ~spriteScaleUpHorizontalReg_21 ? $signed(inSpriteXValue_21) >= 12'sh0 & $signed(
    inSpriteXValue_21) < 12'sh20 : _GEN_1585; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3393 = {{1{spriteYPositionReg_21[9]}},spriteYPositionReg_21}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_21 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3393); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_21 = inSpriteYValue_21[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_21_T = $signed(inSpriteYPreScaled_21) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_21_T_4 = inSpriteYPreScaled_21[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_21_T_8 = _inSpriteVertical_21_T & $signed(inSpriteYPreScaled_21) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_21_T_5 = {$signed(inSpriteYPreScaled_21), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_21_T_14 = _inSpriteVertical_21_T & $signed(inSpriteYPreScaled_21) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1592 = spriteScaleUpVerticalReg_21 ? $signed({{2{_inSpriteY_21_T_4[9]}},_inSpriteY_21_T_4}) :
    $signed(_inSpriteY_21_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1593 = spriteScaleUpVerticalReg_21 ? _inSpriteVertical_21_T_8 : _inSpriteVertical_21_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1594 = ~spriteScaleUpVerticalReg_21 ? $signed({{1{inSpriteYPreScaled_21[10]}},inSpriteYPreScaled_21})
     : $signed(_GEN_1592); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_21 = ~spriteScaleUpVerticalReg_21 ? $signed(inSpriteYPreScaled_21) >= 11'sh0 & $signed(
    inSpriteYPreScaled_21) < 11'sh20 : _GEN_1593; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_22 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_22); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_22_T = $signed(inSpriteXValue_22) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_22_T_4 = inSpriteXValue_22[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_22_T_8 = _inSpriteHorizontal_22_T & $signed(inSpriteXValue_22) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_22_T_5 = {$signed(inSpriteXValue_22), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_22_T_14 = _inSpriteHorizontal_22_T & $signed(inSpriteXValue_22) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1600 = spriteScaleUpHorizontalReg_22 ? $signed({{2{_inSpriteX_22_T_4[10]}},_inSpriteX_22_T_4}) :
    $signed(_inSpriteX_22_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1601 = spriteScaleUpHorizontalReg_22 ? _inSpriteHorizontal_22_T_8 : _inSpriteHorizontal_22_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1602 = ~spriteScaleUpHorizontalReg_22 ? $signed({{1{inSpriteXValue_22[11]}},inSpriteXValue_22}) :
    $signed(_GEN_1600); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_22 = ~spriteScaleUpHorizontalReg_22 ? $signed(inSpriteXValue_22) >= 12'sh0 & $signed(
    inSpriteXValue_22) < 12'sh20 : _GEN_1601; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3395 = {{1{spriteYPositionReg_22[9]}},spriteYPositionReg_22}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_22 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3395); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_22 = inSpriteYValue_22[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_22_T = $signed(inSpriteYPreScaled_22) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_22_T_4 = inSpriteYPreScaled_22[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_22_T_8 = _inSpriteVertical_22_T & $signed(inSpriteYPreScaled_22) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_22_T_5 = {$signed(inSpriteYPreScaled_22), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_22_T_14 = _inSpriteVertical_22_T & $signed(inSpriteYPreScaled_22) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1608 = spriteScaleUpVerticalReg_22 ? $signed({{2{_inSpriteY_22_T_4[9]}},_inSpriteY_22_T_4}) :
    $signed(_inSpriteY_22_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1609 = spriteScaleUpVerticalReg_22 ? _inSpriteVertical_22_T_8 : _inSpriteVertical_22_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1610 = ~spriteScaleUpVerticalReg_22 ? $signed({{1{inSpriteYPreScaled_22[10]}},inSpriteYPreScaled_22})
     : $signed(_GEN_1608); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_22 = ~spriteScaleUpVerticalReg_22 ? $signed(inSpriteYPreScaled_22) >= 11'sh0 & $signed(
    inSpriteYPreScaled_22) < 11'sh20 : _GEN_1609; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_23 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_23); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_23_T = $signed(inSpriteXValue_23) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_23_T_4 = inSpriteXValue_23[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_23_T_8 = _inSpriteHorizontal_23_T & $signed(inSpriteXValue_23) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_23_T_5 = {$signed(inSpriteXValue_23), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_23_T_14 = _inSpriteHorizontal_23_T & $signed(inSpriteXValue_23) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1616 = spriteScaleUpHorizontalReg_23 ? $signed({{2{_inSpriteX_23_T_4[10]}},_inSpriteX_23_T_4}) :
    $signed(_inSpriteX_23_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1617 = spriteScaleUpHorizontalReg_23 ? _inSpriteHorizontal_23_T_8 : _inSpriteHorizontal_23_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1618 = ~spriteScaleUpHorizontalReg_23 ? $signed({{1{inSpriteXValue_23[11]}},inSpriteXValue_23}) :
    $signed(_GEN_1616); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_23 = ~spriteScaleUpHorizontalReg_23 ? $signed(inSpriteXValue_23) >= 12'sh0 & $signed(
    inSpriteXValue_23) < 12'sh20 : _GEN_1617; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3397 = {{1{spriteYPositionReg_23[9]}},spriteYPositionReg_23}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_23 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3397); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_23 = inSpriteYValue_23[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_23_T = $signed(inSpriteYPreScaled_23) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_23_T_4 = inSpriteYPreScaled_23[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_23_T_8 = _inSpriteVertical_23_T & $signed(inSpriteYPreScaled_23) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_23_T_5 = {$signed(inSpriteYPreScaled_23), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_23_T_14 = _inSpriteVertical_23_T & $signed(inSpriteYPreScaled_23) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1624 = spriteScaleUpVerticalReg_23 ? $signed({{2{_inSpriteY_23_T_4[9]}},_inSpriteY_23_T_4}) :
    $signed(_inSpriteY_23_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1625 = spriteScaleUpVerticalReg_23 ? _inSpriteVertical_23_T_8 : _inSpriteVertical_23_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1626 = ~spriteScaleUpVerticalReg_23 ? $signed({{1{inSpriteYPreScaled_23[10]}},inSpriteYPreScaled_23})
     : $signed(_GEN_1624); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_23 = ~spriteScaleUpVerticalReg_23 ? $signed(inSpriteYPreScaled_23) >= 11'sh0 & $signed(
    inSpriteYPreScaled_23) < 11'sh20 : _GEN_1625; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_24 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_24); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_24_T = $signed(inSpriteXValue_24) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_24_T_4 = inSpriteXValue_24[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_24_T_8 = _inSpriteHorizontal_24_T & $signed(inSpriteXValue_24) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_24_T_5 = {$signed(inSpriteXValue_24), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_24_T_14 = _inSpriteHorizontal_24_T & $signed(inSpriteXValue_24) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1632 = spriteScaleUpHorizontalReg_24 ? $signed({{2{_inSpriteX_24_T_4[10]}},_inSpriteX_24_T_4}) :
    $signed(_inSpriteX_24_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1633 = spriteScaleUpHorizontalReg_24 ? _inSpriteHorizontal_24_T_8 : _inSpriteHorizontal_24_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1634 = ~spriteScaleUpHorizontalReg_24 ? $signed({{1{inSpriteXValue_24[11]}},inSpriteXValue_24}) :
    $signed(_GEN_1632); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_24 = ~spriteScaleUpHorizontalReg_24 ? $signed(inSpriteXValue_24) >= 12'sh0 & $signed(
    inSpriteXValue_24) < 12'sh20 : _GEN_1633; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3399 = {{1{spriteYPositionReg_24[9]}},spriteYPositionReg_24}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_24 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3399); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_24 = inSpriteYValue_24[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_24_T = $signed(inSpriteYPreScaled_24) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_24_T_4 = inSpriteYPreScaled_24[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_24_T_8 = _inSpriteVertical_24_T & $signed(inSpriteYPreScaled_24) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_24_T_5 = {$signed(inSpriteYPreScaled_24), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_24_T_14 = _inSpriteVertical_24_T & $signed(inSpriteYPreScaled_24) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1640 = spriteScaleUpVerticalReg_24 ? $signed({{2{_inSpriteY_24_T_4[9]}},_inSpriteY_24_T_4}) :
    $signed(_inSpriteY_24_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1641 = spriteScaleUpVerticalReg_24 ? _inSpriteVertical_24_T_8 : _inSpriteVertical_24_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1642 = ~spriteScaleUpVerticalReg_24 ? $signed({{1{inSpriteYPreScaled_24[10]}},inSpriteYPreScaled_24})
     : $signed(_GEN_1640); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_24 = ~spriteScaleUpVerticalReg_24 ? $signed(inSpriteYPreScaled_24) >= 11'sh0 & $signed(
    inSpriteYPreScaled_24) < 11'sh20 : _GEN_1641; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_25 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_25); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_25_T = $signed(inSpriteXValue_25) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_25_T_4 = inSpriteXValue_25[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_25_T_8 = _inSpriteHorizontal_25_T & $signed(inSpriteXValue_25) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_25_T_5 = {$signed(inSpriteXValue_25), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_25_T_14 = _inSpriteHorizontal_25_T & $signed(inSpriteXValue_25) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1648 = spriteScaleUpHorizontalReg_25 ? $signed({{2{_inSpriteX_25_T_4[10]}},_inSpriteX_25_T_4}) :
    $signed(_inSpriteX_25_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1649 = spriteScaleUpHorizontalReg_25 ? _inSpriteHorizontal_25_T_8 : _inSpriteHorizontal_25_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1650 = ~spriteScaleUpHorizontalReg_25 ? $signed({{1{inSpriteXValue_25[11]}},inSpriteXValue_25}) :
    $signed(_GEN_1648); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_25 = ~spriteScaleUpHorizontalReg_25 ? $signed(inSpriteXValue_25) >= 12'sh0 & $signed(
    inSpriteXValue_25) < 12'sh20 : _GEN_1649; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3401 = {{1{spriteYPositionReg_25[9]}},spriteYPositionReg_25}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_25 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3401); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_25 = inSpriteYValue_25[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_25_T = $signed(inSpriteYPreScaled_25) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_25_T_4 = inSpriteYPreScaled_25[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_25_T_8 = _inSpriteVertical_25_T & $signed(inSpriteYPreScaled_25) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_25_T_5 = {$signed(inSpriteYPreScaled_25), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_25_T_14 = _inSpriteVertical_25_T & $signed(inSpriteYPreScaled_25) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1656 = spriteScaleUpVerticalReg_25 ? $signed({{2{_inSpriteY_25_T_4[9]}},_inSpriteY_25_T_4}) :
    $signed(_inSpriteY_25_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1657 = spriteScaleUpVerticalReg_25 ? _inSpriteVertical_25_T_8 : _inSpriteVertical_25_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1658 = ~spriteScaleUpVerticalReg_25 ? $signed({{1{inSpriteYPreScaled_25[10]}},inSpriteYPreScaled_25})
     : $signed(_GEN_1656); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_25 = ~spriteScaleUpVerticalReg_25 ? $signed(inSpriteYPreScaled_25) >= 11'sh0 & $signed(
    inSpriteYPreScaled_25) < 11'sh20 : _GEN_1657; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_26 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_26); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_26_T = $signed(inSpriteXValue_26) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_26_T_4 = inSpriteXValue_26[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_26_T_8 = _inSpriteHorizontal_26_T & $signed(inSpriteXValue_26) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_26_T_5 = {$signed(inSpriteXValue_26), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_26_T_14 = _inSpriteHorizontal_26_T & $signed(inSpriteXValue_26) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1664 = spriteScaleUpHorizontalReg_26 ? $signed({{2{_inSpriteX_26_T_4[10]}},_inSpriteX_26_T_4}) :
    $signed(_inSpriteX_26_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1665 = spriteScaleUpHorizontalReg_26 ? _inSpriteHorizontal_26_T_8 : _inSpriteHorizontal_26_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1666 = ~spriteScaleUpHorizontalReg_26 ? $signed({{1{inSpriteXValue_26[11]}},inSpriteXValue_26}) :
    $signed(_GEN_1664); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_26 = ~spriteScaleUpHorizontalReg_26 ? $signed(inSpriteXValue_26) >= 12'sh0 & $signed(
    inSpriteXValue_26) < 12'sh20 : _GEN_1665; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3403 = {{1{spriteYPositionReg_26[9]}},spriteYPositionReg_26}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_26 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3403); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_26 = inSpriteYValue_26[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_26_T = $signed(inSpriteYPreScaled_26) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_26_T_4 = inSpriteYPreScaled_26[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_26_T_8 = _inSpriteVertical_26_T & $signed(inSpriteYPreScaled_26) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_26_T_5 = {$signed(inSpriteYPreScaled_26), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_26_T_14 = _inSpriteVertical_26_T & $signed(inSpriteYPreScaled_26) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1672 = spriteScaleUpVerticalReg_26 ? $signed({{2{_inSpriteY_26_T_4[9]}},_inSpriteY_26_T_4}) :
    $signed(_inSpriteY_26_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1673 = spriteScaleUpVerticalReg_26 ? _inSpriteVertical_26_T_8 : _inSpriteVertical_26_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1674 = ~spriteScaleUpVerticalReg_26 ? $signed({{1{inSpriteYPreScaled_26[10]}},inSpriteYPreScaled_26})
     : $signed(_GEN_1672); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_26 = ~spriteScaleUpVerticalReg_26 ? $signed(inSpriteYPreScaled_26) >= 11'sh0 & $signed(
    inSpriteYPreScaled_26) < 11'sh20 : _GEN_1673; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_27 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_27); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_27_T = $signed(inSpriteXValue_27) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_27_T_4 = inSpriteXValue_27[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_27_T_8 = _inSpriteHorizontal_27_T & $signed(inSpriteXValue_27) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_27_T_5 = {$signed(inSpriteXValue_27), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_27_T_14 = _inSpriteHorizontal_27_T & $signed(inSpriteXValue_27) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1680 = spriteScaleUpHorizontalReg_27 ? $signed({{2{_inSpriteX_27_T_4[10]}},_inSpriteX_27_T_4}) :
    $signed(_inSpriteX_27_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1681 = spriteScaleUpHorizontalReg_27 ? _inSpriteHorizontal_27_T_8 : _inSpriteHorizontal_27_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1682 = ~spriteScaleUpHorizontalReg_27 ? $signed({{1{inSpriteXValue_27[11]}},inSpriteXValue_27}) :
    $signed(_GEN_1680); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_27 = ~spriteScaleUpHorizontalReg_27 ? $signed(inSpriteXValue_27) >= 12'sh0 & $signed(
    inSpriteXValue_27) < 12'sh20 : _GEN_1681; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3405 = {{1{spriteYPositionReg_27[9]}},spriteYPositionReg_27}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_27 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3405); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_27 = inSpriteYValue_27[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_27_T = $signed(inSpriteYPreScaled_27) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_27_T_4 = inSpriteYPreScaled_27[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_27_T_8 = _inSpriteVertical_27_T & $signed(inSpriteYPreScaled_27) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_27_T_5 = {$signed(inSpriteYPreScaled_27), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_27_T_14 = _inSpriteVertical_27_T & $signed(inSpriteYPreScaled_27) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1688 = spriteScaleUpVerticalReg_27 ? $signed({{2{_inSpriteY_27_T_4[9]}},_inSpriteY_27_T_4}) :
    $signed(_inSpriteY_27_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1689 = spriteScaleUpVerticalReg_27 ? _inSpriteVertical_27_T_8 : _inSpriteVertical_27_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1690 = ~spriteScaleUpVerticalReg_27 ? $signed({{1{inSpriteYPreScaled_27[10]}},inSpriteYPreScaled_27})
     : $signed(_GEN_1688); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_27 = ~spriteScaleUpVerticalReg_27 ? $signed(inSpriteYPreScaled_27) >= 11'sh0 & $signed(
    inSpriteYPreScaled_27) < 11'sh20 : _GEN_1689; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_28 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_28); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_28_T = $signed(inSpriteXValue_28) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_28_T_4 = inSpriteXValue_28[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_28_T_8 = _inSpriteHorizontal_28_T & $signed(inSpriteXValue_28) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_28_T_5 = {$signed(inSpriteXValue_28), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_28_T_14 = _inSpriteHorizontal_28_T & $signed(inSpriteXValue_28) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1696 = spriteScaleUpHorizontalReg_28 ? $signed({{2{_inSpriteX_28_T_4[10]}},_inSpriteX_28_T_4}) :
    $signed(_inSpriteX_28_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1697 = spriteScaleUpHorizontalReg_28 ? _inSpriteHorizontal_28_T_8 : _inSpriteHorizontal_28_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1698 = ~spriteScaleUpHorizontalReg_28 ? $signed({{1{inSpriteXValue_28[11]}},inSpriteXValue_28}) :
    $signed(_GEN_1696); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_28 = ~spriteScaleUpHorizontalReg_28 ? $signed(inSpriteXValue_28) >= 12'sh0 & $signed(
    inSpriteXValue_28) < 12'sh20 : _GEN_1697; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3407 = {{1{spriteYPositionReg_28[9]}},spriteYPositionReg_28}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_28 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3407); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_28 = inSpriteYValue_28[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_28_T = $signed(inSpriteYPreScaled_28) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_28_T_4 = inSpriteYPreScaled_28[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_28_T_8 = _inSpriteVertical_28_T & $signed(inSpriteYPreScaled_28) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_28_T_5 = {$signed(inSpriteYPreScaled_28), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_28_T_14 = _inSpriteVertical_28_T & $signed(inSpriteYPreScaled_28) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1704 = spriteScaleUpVerticalReg_28 ? $signed({{2{_inSpriteY_28_T_4[9]}},_inSpriteY_28_T_4}) :
    $signed(_inSpriteY_28_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1705 = spriteScaleUpVerticalReg_28 ? _inSpriteVertical_28_T_8 : _inSpriteVertical_28_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1706 = ~spriteScaleUpVerticalReg_28 ? $signed({{1{inSpriteYPreScaled_28[10]}},inSpriteYPreScaled_28})
     : $signed(_GEN_1704); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_28 = ~spriteScaleUpVerticalReg_28 ? $signed(inSpriteYPreScaled_28) >= 11'sh0 & $signed(
    inSpriteYPreScaled_28) < 11'sh20 : _GEN_1705; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_29 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_29); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_29_T = $signed(inSpriteXValue_29) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_29_T_4 = inSpriteXValue_29[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_29_T_8 = _inSpriteHorizontal_29_T & $signed(inSpriteXValue_29) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_29_T_5 = {$signed(inSpriteXValue_29), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_29_T_14 = _inSpriteHorizontal_29_T & $signed(inSpriteXValue_29) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1712 = spriteScaleUpHorizontalReg_29 ? $signed({{2{_inSpriteX_29_T_4[10]}},_inSpriteX_29_T_4}) :
    $signed(_inSpriteX_29_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1713 = spriteScaleUpHorizontalReg_29 ? _inSpriteHorizontal_29_T_8 : _inSpriteHorizontal_29_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1714 = ~spriteScaleUpHorizontalReg_29 ? $signed({{1{inSpriteXValue_29[11]}},inSpriteXValue_29}) :
    $signed(_GEN_1712); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_29 = ~spriteScaleUpHorizontalReg_29 ? $signed(inSpriteXValue_29) >= 12'sh0 & $signed(
    inSpriteXValue_29) < 12'sh20 : _GEN_1713; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3409 = {{1{spriteYPositionReg_29[9]}},spriteYPositionReg_29}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_29 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3409); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_29 = inSpriteYValue_29[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_29_T = $signed(inSpriteYPreScaled_29) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_29_T_4 = inSpriteYPreScaled_29[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_29_T_8 = _inSpriteVertical_29_T & $signed(inSpriteYPreScaled_29) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_29_T_5 = {$signed(inSpriteYPreScaled_29), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_29_T_14 = _inSpriteVertical_29_T & $signed(inSpriteYPreScaled_29) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1720 = spriteScaleUpVerticalReg_29 ? $signed({{2{_inSpriteY_29_T_4[9]}},_inSpriteY_29_T_4}) :
    $signed(_inSpriteY_29_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1721 = spriteScaleUpVerticalReg_29 ? _inSpriteVertical_29_T_8 : _inSpriteVertical_29_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1722 = ~spriteScaleUpVerticalReg_29 ? $signed({{1{inSpriteYPreScaled_29[10]}},inSpriteYPreScaled_29})
     : $signed(_GEN_1720); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_29 = ~spriteScaleUpVerticalReg_29 ? $signed(inSpriteYPreScaled_29) >= 11'sh0 & $signed(
    inSpriteYPreScaled_29) < 11'sh20 : _GEN_1721; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_30 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_30); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_30_T = $signed(inSpriteXValue_30) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_30_T_4 = inSpriteXValue_30[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_30_T_8 = _inSpriteHorizontal_30_T & $signed(inSpriteXValue_30) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_30_T_5 = {$signed(inSpriteXValue_30), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_30_T_14 = _inSpriteHorizontal_30_T & $signed(inSpriteXValue_30) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1728 = spriteScaleUpHorizontalReg_30 ? $signed({{2{_inSpriteX_30_T_4[10]}},_inSpriteX_30_T_4}) :
    $signed(_inSpriteX_30_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1729 = spriteScaleUpHorizontalReg_30 ? _inSpriteHorizontal_30_T_8 : _inSpriteHorizontal_30_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1730 = ~spriteScaleUpHorizontalReg_30 ? $signed({{1{inSpriteXValue_30[11]}},inSpriteXValue_30}) :
    $signed(_GEN_1728); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_30 = ~spriteScaleUpHorizontalReg_30 ? $signed(inSpriteXValue_30) >= 12'sh0 & $signed(
    inSpriteXValue_30) < 12'sh20 : _GEN_1729; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3411 = {{1{spriteYPositionReg_30[9]}},spriteYPositionReg_30}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_30 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3411); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_30 = inSpriteYValue_30[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_30_T = $signed(inSpriteYPreScaled_30) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_30_T_4 = inSpriteYPreScaled_30[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_30_T_8 = _inSpriteVertical_30_T & $signed(inSpriteYPreScaled_30) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_30_T_5 = {$signed(inSpriteYPreScaled_30), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_30_T_14 = _inSpriteVertical_30_T & $signed(inSpriteYPreScaled_30) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1736 = spriteScaleUpVerticalReg_30 ? $signed({{2{_inSpriteY_30_T_4[9]}},_inSpriteY_30_T_4}) :
    $signed(_inSpriteY_30_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1737 = spriteScaleUpVerticalReg_30 ? _inSpriteVertical_30_T_8 : _inSpriteVertical_30_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1738 = ~spriteScaleUpVerticalReg_30 ? $signed({{1{inSpriteYPreScaled_30[10]}},inSpriteYPreScaled_30})
     : $signed(_GEN_1736); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_30 = ~spriteScaleUpVerticalReg_30 ? $signed(inSpriteYPreScaled_30) >= 11'sh0 & $signed(
    inSpriteYPreScaled_30) < 11'sh20 : _GEN_1737; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_31 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_31); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_31_T = $signed(inSpriteXValue_31) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_31_T_4 = inSpriteXValue_31[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_31_T_8 = _inSpriteHorizontal_31_T & $signed(inSpriteXValue_31) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_31_T_5 = {$signed(inSpriteXValue_31), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_31_T_14 = _inSpriteHorizontal_31_T & $signed(inSpriteXValue_31) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1744 = spriteScaleUpHorizontalReg_31 ? $signed({{2{_inSpriteX_31_T_4[10]}},_inSpriteX_31_T_4}) :
    $signed(_inSpriteX_31_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1745 = spriteScaleUpHorizontalReg_31 ? _inSpriteHorizontal_31_T_8 : _inSpriteHorizontal_31_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1746 = ~spriteScaleUpHorizontalReg_31 ? $signed({{1{inSpriteXValue_31[11]}},inSpriteXValue_31}) :
    $signed(_GEN_1744); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_31 = ~spriteScaleUpHorizontalReg_31 ? $signed(inSpriteXValue_31) >= 12'sh0 & $signed(
    inSpriteXValue_31) < 12'sh20 : _GEN_1745; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3413 = {{1{spriteYPositionReg_31[9]}},spriteYPositionReg_31}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_31 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3413); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_31 = inSpriteYValue_31[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_31_T = $signed(inSpriteYPreScaled_31) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_31_T_4 = inSpriteYPreScaled_31[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_31_T_8 = _inSpriteVertical_31_T & $signed(inSpriteYPreScaled_31) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_31_T_5 = {$signed(inSpriteYPreScaled_31), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_31_T_14 = _inSpriteVertical_31_T & $signed(inSpriteYPreScaled_31) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1752 = spriteScaleUpVerticalReg_31 ? $signed({{2{_inSpriteY_31_T_4[9]}},_inSpriteY_31_T_4}) :
    $signed(_inSpriteY_31_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1753 = spriteScaleUpVerticalReg_31 ? _inSpriteVertical_31_T_8 : _inSpriteVertical_31_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1754 = ~spriteScaleUpVerticalReg_31 ? $signed({{1{inSpriteYPreScaled_31[10]}},inSpriteYPreScaled_31})
     : $signed(_GEN_1752); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_31 = ~spriteScaleUpVerticalReg_31 ? $signed(inSpriteYPreScaled_31) >= 11'sh0 & $signed(
    inSpriteYPreScaled_31) < 11'sh20 : _GEN_1753; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_32 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_32); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_32_T = $signed(inSpriteXValue_32) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_32_T_4 = inSpriteXValue_32[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_32_T_8 = _inSpriteHorizontal_32_T & $signed(inSpriteXValue_32) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_32_T_5 = {$signed(inSpriteXValue_32), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_32_T_14 = _inSpriteHorizontal_32_T & $signed(inSpriteXValue_32) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1760 = spriteScaleUpHorizontalReg_32 ? $signed({{2{_inSpriteX_32_T_4[10]}},_inSpriteX_32_T_4}) :
    $signed(_inSpriteX_32_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1761 = spriteScaleUpHorizontalReg_32 ? _inSpriteHorizontal_32_T_8 : _inSpriteHorizontal_32_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1762 = ~spriteScaleUpHorizontalReg_32 ? $signed({{1{inSpriteXValue_32[11]}},inSpriteXValue_32}) :
    $signed(_GEN_1760); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_32 = ~spriteScaleUpHorizontalReg_32 ? $signed(inSpriteXValue_32) >= 12'sh0 & $signed(
    inSpriteXValue_32) < 12'sh20 : _GEN_1761; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3415 = {{1{spriteYPositionReg_32[9]}},spriteYPositionReg_32}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_32 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3415); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_32 = inSpriteYValue_32[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_32_T = $signed(inSpriteYPreScaled_32) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_32_T_4 = inSpriteYPreScaled_32[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_32_T_8 = _inSpriteVertical_32_T & $signed(inSpriteYPreScaled_32) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_32_T_5 = {$signed(inSpriteYPreScaled_32), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_32_T_14 = _inSpriteVertical_32_T & $signed(inSpriteYPreScaled_32) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1768 = spriteScaleUpVerticalReg_32 ? $signed({{2{_inSpriteY_32_T_4[9]}},_inSpriteY_32_T_4}) :
    $signed(_inSpriteY_32_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1769 = spriteScaleUpVerticalReg_32 ? _inSpriteVertical_32_T_8 : _inSpriteVertical_32_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1770 = ~spriteScaleUpVerticalReg_32 ? $signed({{1{inSpriteYPreScaled_32[10]}},inSpriteYPreScaled_32})
     : $signed(_GEN_1768); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_32 = ~spriteScaleUpVerticalReg_32 ? $signed(inSpriteYPreScaled_32) >= 11'sh0 & $signed(
    inSpriteYPreScaled_32) < 11'sh20 : _GEN_1769; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_33 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_33); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_33_T = $signed(inSpriteXValue_33) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_33_T_4 = inSpriteXValue_33[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_33_T_8 = _inSpriteHorizontal_33_T & $signed(inSpriteXValue_33) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_33_T_5 = {$signed(inSpriteXValue_33), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_33_T_14 = _inSpriteHorizontal_33_T & $signed(inSpriteXValue_33) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1776 = spriteScaleUpHorizontalReg_33 ? $signed({{2{_inSpriteX_33_T_4[10]}},_inSpriteX_33_T_4}) :
    $signed(_inSpriteX_33_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1777 = spriteScaleUpHorizontalReg_33 ? _inSpriteHorizontal_33_T_8 : _inSpriteHorizontal_33_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1778 = ~spriteScaleUpHorizontalReg_33 ? $signed({{1{inSpriteXValue_33[11]}},inSpriteXValue_33}) :
    $signed(_GEN_1776); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_33 = ~spriteScaleUpHorizontalReg_33 ? $signed(inSpriteXValue_33) >= 12'sh0 & $signed(
    inSpriteXValue_33) < 12'sh20 : _GEN_1777; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3417 = {{1{spriteYPositionReg_33[9]}},spriteYPositionReg_33}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_33 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3417); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_33 = inSpriteYValue_33[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_33_T = $signed(inSpriteYPreScaled_33) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_33_T_4 = inSpriteYPreScaled_33[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_33_T_8 = _inSpriteVertical_33_T & $signed(inSpriteYPreScaled_33) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_33_T_5 = {$signed(inSpriteYPreScaled_33), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_33_T_14 = _inSpriteVertical_33_T & $signed(inSpriteYPreScaled_33) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1784 = spriteScaleUpVerticalReg_33 ? $signed({{2{_inSpriteY_33_T_4[9]}},_inSpriteY_33_T_4}) :
    $signed(_inSpriteY_33_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1785 = spriteScaleUpVerticalReg_33 ? _inSpriteVertical_33_T_8 : _inSpriteVertical_33_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1786 = ~spriteScaleUpVerticalReg_33 ? $signed({{1{inSpriteYPreScaled_33[10]}},inSpriteYPreScaled_33})
     : $signed(_GEN_1784); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_33 = ~spriteScaleUpVerticalReg_33 ? $signed(inSpriteYPreScaled_33) >= 11'sh0 & $signed(
    inSpriteYPreScaled_33) < 11'sh20 : _GEN_1785; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_34 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_34); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_34_T = $signed(inSpriteXValue_34) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_34_T_4 = inSpriteXValue_34[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_34_T_8 = _inSpriteHorizontal_34_T & $signed(inSpriteXValue_34) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_34_T_5 = {$signed(inSpriteXValue_34), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_34_T_14 = _inSpriteHorizontal_34_T & $signed(inSpriteXValue_34) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1792 = spriteScaleUpHorizontalReg_34 ? $signed({{2{_inSpriteX_34_T_4[10]}},_inSpriteX_34_T_4}) :
    $signed(_inSpriteX_34_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1793 = spriteScaleUpHorizontalReg_34 ? _inSpriteHorizontal_34_T_8 : _inSpriteHorizontal_34_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1794 = ~spriteScaleUpHorizontalReg_34 ? $signed({{1{inSpriteXValue_34[11]}},inSpriteXValue_34}) :
    $signed(_GEN_1792); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_34 = ~spriteScaleUpHorizontalReg_34 ? $signed(inSpriteXValue_34) >= 12'sh0 & $signed(
    inSpriteXValue_34) < 12'sh20 : _GEN_1793; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3419 = {{1{spriteYPositionReg_34[9]}},spriteYPositionReg_34}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_34 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3419); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_34 = inSpriteYValue_34[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_34_T = $signed(inSpriteYPreScaled_34) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_34_T_4 = inSpriteYPreScaled_34[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_34_T_8 = _inSpriteVertical_34_T & $signed(inSpriteYPreScaled_34) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_34_T_5 = {$signed(inSpriteYPreScaled_34), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_34_T_14 = _inSpriteVertical_34_T & $signed(inSpriteYPreScaled_34) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1800 = spriteScaleUpVerticalReg_34 ? $signed({{2{_inSpriteY_34_T_4[9]}},_inSpriteY_34_T_4}) :
    $signed(_inSpriteY_34_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1801 = spriteScaleUpVerticalReg_34 ? _inSpriteVertical_34_T_8 : _inSpriteVertical_34_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1802 = ~spriteScaleUpVerticalReg_34 ? $signed({{1{inSpriteYPreScaled_34[10]}},inSpriteYPreScaled_34})
     : $signed(_GEN_1800); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_34 = ~spriteScaleUpVerticalReg_34 ? $signed(inSpriteYPreScaled_34) >= 11'sh0 & $signed(
    inSpriteYPreScaled_34) < 11'sh20 : _GEN_1801; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_35 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_35); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_35_T = $signed(inSpriteXValue_35) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_35_T_4 = inSpriteXValue_35[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_35_T_8 = _inSpriteHorizontal_35_T & $signed(inSpriteXValue_35) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_35_T_5 = {$signed(inSpriteXValue_35), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_35_T_14 = _inSpriteHorizontal_35_T & $signed(inSpriteXValue_35) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1808 = spriteScaleUpHorizontalReg_35 ? $signed({{2{_inSpriteX_35_T_4[10]}},_inSpriteX_35_T_4}) :
    $signed(_inSpriteX_35_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1809 = spriteScaleUpHorizontalReg_35 ? _inSpriteHorizontal_35_T_8 : _inSpriteHorizontal_35_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1810 = ~spriteScaleUpHorizontalReg_35 ? $signed({{1{inSpriteXValue_35[11]}},inSpriteXValue_35}) :
    $signed(_GEN_1808); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_35 = ~spriteScaleUpHorizontalReg_35 ? $signed(inSpriteXValue_35) >= 12'sh0 & $signed(
    inSpriteXValue_35) < 12'sh20 : _GEN_1809; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3421 = {{1{spriteYPositionReg_35[9]}},spriteYPositionReg_35}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_35 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3421); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_35 = inSpriteYValue_35[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_35_T = $signed(inSpriteYPreScaled_35) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_35_T_4 = inSpriteYPreScaled_35[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_35_T_8 = _inSpriteVertical_35_T & $signed(inSpriteYPreScaled_35) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_35_T_5 = {$signed(inSpriteYPreScaled_35), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_35_T_14 = _inSpriteVertical_35_T & $signed(inSpriteYPreScaled_35) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1816 = spriteScaleUpVerticalReg_35 ? $signed({{2{_inSpriteY_35_T_4[9]}},_inSpriteY_35_T_4}) :
    $signed(_inSpriteY_35_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1817 = spriteScaleUpVerticalReg_35 ? _inSpriteVertical_35_T_8 : _inSpriteVertical_35_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1818 = ~spriteScaleUpVerticalReg_35 ? $signed({{1{inSpriteYPreScaled_35[10]}},inSpriteYPreScaled_35})
     : $signed(_GEN_1816); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_35 = ~spriteScaleUpVerticalReg_35 ? $signed(inSpriteYPreScaled_35) >= 11'sh0 & $signed(
    inSpriteYPreScaled_35) < 11'sh20 : _GEN_1817; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_36 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_36); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_36_T = $signed(inSpriteXValue_36) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_36_T_4 = inSpriteXValue_36[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_36_T_8 = _inSpriteHorizontal_36_T & $signed(inSpriteXValue_36) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_36_T_5 = {$signed(inSpriteXValue_36), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_36_T_14 = _inSpriteHorizontal_36_T & $signed(inSpriteXValue_36) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1824 = spriteScaleUpHorizontalReg_36 ? $signed({{2{_inSpriteX_36_T_4[10]}},_inSpriteX_36_T_4}) :
    $signed(_inSpriteX_36_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1825 = spriteScaleUpHorizontalReg_36 ? _inSpriteHorizontal_36_T_8 : _inSpriteHorizontal_36_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1826 = ~spriteScaleUpHorizontalReg_36 ? $signed({{1{inSpriteXValue_36[11]}},inSpriteXValue_36}) :
    $signed(_GEN_1824); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_36 = ~spriteScaleUpHorizontalReg_36 ? $signed(inSpriteXValue_36) >= 12'sh0 & $signed(
    inSpriteXValue_36) < 12'sh20 : _GEN_1825; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3423 = {{1{spriteYPositionReg_36[9]}},spriteYPositionReg_36}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_36 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3423); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_36 = inSpriteYValue_36[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_36_T = $signed(inSpriteYPreScaled_36) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_36_T_4 = inSpriteYPreScaled_36[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_36_T_8 = _inSpriteVertical_36_T & $signed(inSpriteYPreScaled_36) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_36_T_5 = {$signed(inSpriteYPreScaled_36), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_36_T_14 = _inSpriteVertical_36_T & $signed(inSpriteYPreScaled_36) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1832 = spriteScaleUpVerticalReg_36 ? $signed({{2{_inSpriteY_36_T_4[9]}},_inSpriteY_36_T_4}) :
    $signed(_inSpriteY_36_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1833 = spriteScaleUpVerticalReg_36 ? _inSpriteVertical_36_T_8 : _inSpriteVertical_36_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1834 = ~spriteScaleUpVerticalReg_36 ? $signed({{1{inSpriteYPreScaled_36[10]}},inSpriteYPreScaled_36})
     : $signed(_GEN_1832); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_36 = ~spriteScaleUpVerticalReg_36 ? $signed(inSpriteYPreScaled_36) >= 11'sh0 & $signed(
    inSpriteYPreScaled_36) < 11'sh20 : _GEN_1833; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_37 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_37); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_37_T = $signed(inSpriteXValue_37) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_37_T_4 = inSpriteXValue_37[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_37_T_8 = _inSpriteHorizontal_37_T & $signed(inSpriteXValue_37) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_37_T_5 = {$signed(inSpriteXValue_37), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_37_T_14 = _inSpriteHorizontal_37_T & $signed(inSpriteXValue_37) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1840 = spriteScaleUpHorizontalReg_37 ? $signed({{2{_inSpriteX_37_T_4[10]}},_inSpriteX_37_T_4}) :
    $signed(_inSpriteX_37_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1841 = spriteScaleUpHorizontalReg_37 ? _inSpriteHorizontal_37_T_8 : _inSpriteHorizontal_37_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1842 = ~spriteScaleUpHorizontalReg_37 ? $signed({{1{inSpriteXValue_37[11]}},inSpriteXValue_37}) :
    $signed(_GEN_1840); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_37 = ~spriteScaleUpHorizontalReg_37 ? $signed(inSpriteXValue_37) >= 12'sh0 & $signed(
    inSpriteXValue_37) < 12'sh20 : _GEN_1841; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3425 = {{1{spriteYPositionReg_37[9]}},spriteYPositionReg_37}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_37 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3425); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_37 = inSpriteYValue_37[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_37_T = $signed(inSpriteYPreScaled_37) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_37_T_4 = inSpriteYPreScaled_37[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_37_T_8 = _inSpriteVertical_37_T & $signed(inSpriteYPreScaled_37) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_37_T_5 = {$signed(inSpriteYPreScaled_37), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_37_T_14 = _inSpriteVertical_37_T & $signed(inSpriteYPreScaled_37) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1848 = spriteScaleUpVerticalReg_37 ? $signed({{2{_inSpriteY_37_T_4[9]}},_inSpriteY_37_T_4}) :
    $signed(_inSpriteY_37_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1849 = spriteScaleUpVerticalReg_37 ? _inSpriteVertical_37_T_8 : _inSpriteVertical_37_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1850 = ~spriteScaleUpVerticalReg_37 ? $signed({{1{inSpriteYPreScaled_37[10]}},inSpriteYPreScaled_37})
     : $signed(_GEN_1848); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_37 = ~spriteScaleUpVerticalReg_37 ? $signed(inSpriteYPreScaled_37) >= 11'sh0 & $signed(
    inSpriteYPreScaled_37) < 11'sh20 : _GEN_1849; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_38 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_38); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_38_T = $signed(inSpriteXValue_38) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_38_T_4 = inSpriteXValue_38[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_38_T_8 = _inSpriteHorizontal_38_T & $signed(inSpriteXValue_38) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_38_T_5 = {$signed(inSpriteXValue_38), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_38_T_14 = _inSpriteHorizontal_38_T & $signed(inSpriteXValue_38) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1856 = spriteScaleUpHorizontalReg_38 ? $signed({{2{_inSpriteX_38_T_4[10]}},_inSpriteX_38_T_4}) :
    $signed(_inSpriteX_38_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1857 = spriteScaleUpHorizontalReg_38 ? _inSpriteHorizontal_38_T_8 : _inSpriteHorizontal_38_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1858 = ~spriteScaleUpHorizontalReg_38 ? $signed({{1{inSpriteXValue_38[11]}},inSpriteXValue_38}) :
    $signed(_GEN_1856); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_38 = ~spriteScaleUpHorizontalReg_38 ? $signed(inSpriteXValue_38) >= 12'sh0 & $signed(
    inSpriteXValue_38) < 12'sh20 : _GEN_1857; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3427 = {{1{spriteYPositionReg_38[9]}},spriteYPositionReg_38}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_38 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3427); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_38 = inSpriteYValue_38[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_38_T = $signed(inSpriteYPreScaled_38) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_38_T_4 = inSpriteYPreScaled_38[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_38_T_8 = _inSpriteVertical_38_T & $signed(inSpriteYPreScaled_38) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_38_T_5 = {$signed(inSpriteYPreScaled_38), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_38_T_14 = _inSpriteVertical_38_T & $signed(inSpriteYPreScaled_38) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1864 = spriteScaleUpVerticalReg_38 ? $signed({{2{_inSpriteY_38_T_4[9]}},_inSpriteY_38_T_4}) :
    $signed(_inSpriteY_38_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1865 = spriteScaleUpVerticalReg_38 ? _inSpriteVertical_38_T_8 : _inSpriteVertical_38_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1866 = ~spriteScaleUpVerticalReg_38 ? $signed({{1{inSpriteYPreScaled_38[10]}},inSpriteYPreScaled_38})
     : $signed(_GEN_1864); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_38 = ~spriteScaleUpVerticalReg_38 ? $signed(inSpriteYPreScaled_38) >= 11'sh0 & $signed(
    inSpriteYPreScaled_38) < 11'sh20 : _GEN_1865; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_39 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_39); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_39_T = $signed(inSpriteXValue_39) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_39_T_4 = inSpriteXValue_39[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_39_T_8 = _inSpriteHorizontal_39_T & $signed(inSpriteXValue_39) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_39_T_5 = {$signed(inSpriteXValue_39), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_39_T_14 = _inSpriteHorizontal_39_T & $signed(inSpriteXValue_39) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1872 = spriteScaleUpHorizontalReg_39 ? $signed({{2{_inSpriteX_39_T_4[10]}},_inSpriteX_39_T_4}) :
    $signed(_inSpriteX_39_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1873 = spriteScaleUpHorizontalReg_39 ? _inSpriteHorizontal_39_T_8 : _inSpriteHorizontal_39_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1874 = ~spriteScaleUpHorizontalReg_39 ? $signed({{1{inSpriteXValue_39[11]}},inSpriteXValue_39}) :
    $signed(_GEN_1872); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_39 = ~spriteScaleUpHorizontalReg_39 ? $signed(inSpriteXValue_39) >= 12'sh0 & $signed(
    inSpriteXValue_39) < 12'sh20 : _GEN_1873; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3429 = {{1{spriteYPositionReg_39[9]}},spriteYPositionReg_39}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_39 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3429); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_39 = inSpriteYValue_39[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_39_T = $signed(inSpriteYPreScaled_39) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_39_T_4 = inSpriteYPreScaled_39[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_39_T_8 = _inSpriteVertical_39_T & $signed(inSpriteYPreScaled_39) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_39_T_5 = {$signed(inSpriteYPreScaled_39), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_39_T_14 = _inSpriteVertical_39_T & $signed(inSpriteYPreScaled_39) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1880 = spriteScaleUpVerticalReg_39 ? $signed({{2{_inSpriteY_39_T_4[9]}},_inSpriteY_39_T_4}) :
    $signed(_inSpriteY_39_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1881 = spriteScaleUpVerticalReg_39 ? _inSpriteVertical_39_T_8 : _inSpriteVertical_39_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1882 = ~spriteScaleUpVerticalReg_39 ? $signed({{1{inSpriteYPreScaled_39[10]}},inSpriteYPreScaled_39})
     : $signed(_GEN_1880); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_39 = ~spriteScaleUpVerticalReg_39 ? $signed(inSpriteYPreScaled_39) >= 11'sh0 & $signed(
    inSpriteYPreScaled_39) < 11'sh20 : _GEN_1881; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_40 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_40); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_40_T = $signed(inSpriteXValue_40) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_40_T_4 = inSpriteXValue_40[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_40_T_8 = _inSpriteHorizontal_40_T & $signed(inSpriteXValue_40) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_40_T_5 = {$signed(inSpriteXValue_40), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_40_T_14 = _inSpriteHorizontal_40_T & $signed(inSpriteXValue_40) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1888 = spriteScaleUpHorizontalReg_40 ? $signed({{2{_inSpriteX_40_T_4[10]}},_inSpriteX_40_T_4}) :
    $signed(_inSpriteX_40_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1889 = spriteScaleUpHorizontalReg_40 ? _inSpriteHorizontal_40_T_8 : _inSpriteHorizontal_40_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1890 = ~spriteScaleUpHorizontalReg_40 ? $signed({{1{inSpriteXValue_40[11]}},inSpriteXValue_40}) :
    $signed(_GEN_1888); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_40 = ~spriteScaleUpHorizontalReg_40 ? $signed(inSpriteXValue_40) >= 12'sh0 & $signed(
    inSpriteXValue_40) < 12'sh20 : _GEN_1889; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3431 = {{1{spriteYPositionReg_40[9]}},spriteYPositionReg_40}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_40 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3431); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_40 = inSpriteYValue_40[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_40_T = $signed(inSpriteYPreScaled_40) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_40_T_4 = inSpriteYPreScaled_40[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_40_T_8 = _inSpriteVertical_40_T & $signed(inSpriteYPreScaled_40) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_40_T_5 = {$signed(inSpriteYPreScaled_40), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_40_T_14 = _inSpriteVertical_40_T & $signed(inSpriteYPreScaled_40) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1896 = spriteScaleUpVerticalReg_40 ? $signed({{2{_inSpriteY_40_T_4[9]}},_inSpriteY_40_T_4}) :
    $signed(_inSpriteY_40_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1897 = spriteScaleUpVerticalReg_40 ? _inSpriteVertical_40_T_8 : _inSpriteVertical_40_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1898 = ~spriteScaleUpVerticalReg_40 ? $signed({{1{inSpriteYPreScaled_40[10]}},inSpriteYPreScaled_40})
     : $signed(_GEN_1896); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_40 = ~spriteScaleUpVerticalReg_40 ? $signed(inSpriteYPreScaled_40) >= 11'sh0 & $signed(
    inSpriteYPreScaled_40) < 11'sh20 : _GEN_1897; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_41 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_41); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_41_T = $signed(inSpriteXValue_41) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_41_T_4 = inSpriteXValue_41[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_41_T_8 = _inSpriteHorizontal_41_T & $signed(inSpriteXValue_41) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_41_T_5 = {$signed(inSpriteXValue_41), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_41_T_14 = _inSpriteHorizontal_41_T & $signed(inSpriteXValue_41) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1904 = spriteScaleUpHorizontalReg_41 ? $signed({{2{_inSpriteX_41_T_4[10]}},_inSpriteX_41_T_4}) :
    $signed(_inSpriteX_41_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1905 = spriteScaleUpHorizontalReg_41 ? _inSpriteHorizontal_41_T_8 : _inSpriteHorizontal_41_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1906 = ~spriteScaleUpHorizontalReg_41 ? $signed({{1{inSpriteXValue_41[11]}},inSpriteXValue_41}) :
    $signed(_GEN_1904); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_41 = ~spriteScaleUpHorizontalReg_41 ? $signed(inSpriteXValue_41) >= 12'sh0 & $signed(
    inSpriteXValue_41) < 12'sh20 : _GEN_1905; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3433 = {{1{spriteYPositionReg_41[9]}},spriteYPositionReg_41}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_41 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3433); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_41 = inSpriteYValue_41[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_41_T = $signed(inSpriteYPreScaled_41) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_41_T_4 = inSpriteYPreScaled_41[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_41_T_8 = _inSpriteVertical_41_T & $signed(inSpriteYPreScaled_41) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_41_T_5 = {$signed(inSpriteYPreScaled_41), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_41_T_14 = _inSpriteVertical_41_T & $signed(inSpriteYPreScaled_41) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1912 = spriteScaleUpVerticalReg_41 ? $signed({{2{_inSpriteY_41_T_4[9]}},_inSpriteY_41_T_4}) :
    $signed(_inSpriteY_41_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1913 = spriteScaleUpVerticalReg_41 ? _inSpriteVertical_41_T_8 : _inSpriteVertical_41_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1914 = ~spriteScaleUpVerticalReg_41 ? $signed({{1{inSpriteYPreScaled_41[10]}},inSpriteYPreScaled_41})
     : $signed(_GEN_1912); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_41 = ~spriteScaleUpVerticalReg_41 ? $signed(inSpriteYPreScaled_41) >= 11'sh0 & $signed(
    inSpriteYPreScaled_41) < 11'sh20 : _GEN_1913; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_42 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_42); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_42_T = $signed(inSpriteXValue_42) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_42_T_4 = inSpriteXValue_42[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_42_T_8 = _inSpriteHorizontal_42_T & $signed(inSpriteXValue_42) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_42_T_5 = {$signed(inSpriteXValue_42), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_42_T_14 = _inSpriteHorizontal_42_T & $signed(inSpriteXValue_42) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1920 = spriteScaleUpHorizontalReg_42 ? $signed({{2{_inSpriteX_42_T_4[10]}},_inSpriteX_42_T_4}) :
    $signed(_inSpriteX_42_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1921 = spriteScaleUpHorizontalReg_42 ? _inSpriteHorizontal_42_T_8 : _inSpriteHorizontal_42_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1922 = ~spriteScaleUpHorizontalReg_42 ? $signed({{1{inSpriteXValue_42[11]}},inSpriteXValue_42}) :
    $signed(_GEN_1920); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_42 = ~spriteScaleUpHorizontalReg_42 ? $signed(inSpriteXValue_42) >= 12'sh0 & $signed(
    inSpriteXValue_42) < 12'sh20 : _GEN_1921; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3435 = {{1{spriteYPositionReg_42[9]}},spriteYPositionReg_42}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_42 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3435); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_42 = inSpriteYValue_42[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_42_T = $signed(inSpriteYPreScaled_42) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_42_T_4 = inSpriteYPreScaled_42[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_42_T_8 = _inSpriteVertical_42_T & $signed(inSpriteYPreScaled_42) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_42_T_5 = {$signed(inSpriteYPreScaled_42), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_42_T_14 = _inSpriteVertical_42_T & $signed(inSpriteYPreScaled_42) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1928 = spriteScaleUpVerticalReg_42 ? $signed({{2{_inSpriteY_42_T_4[9]}},_inSpriteY_42_T_4}) :
    $signed(_inSpriteY_42_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1929 = spriteScaleUpVerticalReg_42 ? _inSpriteVertical_42_T_8 : _inSpriteVertical_42_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1930 = ~spriteScaleUpVerticalReg_42 ? $signed({{1{inSpriteYPreScaled_42[10]}},inSpriteYPreScaled_42})
     : $signed(_GEN_1928); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_42 = ~spriteScaleUpVerticalReg_42 ? $signed(inSpriteYPreScaled_42) >= 11'sh0 & $signed(
    inSpriteYPreScaled_42) < 11'sh20 : _GEN_1929; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_43 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_43); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_43_T = $signed(inSpriteXValue_43) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_43_T_4 = inSpriteXValue_43[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_43_T_8 = _inSpriteHorizontal_43_T & $signed(inSpriteXValue_43) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_43_T_5 = {$signed(inSpriteXValue_43), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_43_T_14 = _inSpriteHorizontal_43_T & $signed(inSpriteXValue_43) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1936 = spriteScaleUpHorizontalReg_43 ? $signed({{2{_inSpriteX_43_T_4[10]}},_inSpriteX_43_T_4}) :
    $signed(_inSpriteX_43_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1937 = spriteScaleUpHorizontalReg_43 ? _inSpriteHorizontal_43_T_8 : _inSpriteHorizontal_43_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1938 = ~spriteScaleUpHorizontalReg_43 ? $signed({{1{inSpriteXValue_43[11]}},inSpriteXValue_43}) :
    $signed(_GEN_1936); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_43 = ~spriteScaleUpHorizontalReg_43 ? $signed(inSpriteXValue_43) >= 12'sh0 & $signed(
    inSpriteXValue_43) < 12'sh20 : _GEN_1937; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3437 = {{1{spriteYPositionReg_43[9]}},spriteYPositionReg_43}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_43 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3437); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_43 = inSpriteYValue_43[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_43_T = $signed(inSpriteYPreScaled_43) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_43_T_4 = inSpriteYPreScaled_43[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_43_T_8 = _inSpriteVertical_43_T & $signed(inSpriteYPreScaled_43) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_43_T_5 = {$signed(inSpriteYPreScaled_43), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_43_T_14 = _inSpriteVertical_43_T & $signed(inSpriteYPreScaled_43) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1944 = spriteScaleUpVerticalReg_43 ? $signed({{2{_inSpriteY_43_T_4[9]}},_inSpriteY_43_T_4}) :
    $signed(_inSpriteY_43_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1945 = spriteScaleUpVerticalReg_43 ? _inSpriteVertical_43_T_8 : _inSpriteVertical_43_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1946 = ~spriteScaleUpVerticalReg_43 ? $signed({{1{inSpriteYPreScaled_43[10]}},inSpriteYPreScaled_43})
     : $signed(_GEN_1944); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_43 = ~spriteScaleUpVerticalReg_43 ? $signed(inSpriteYPreScaled_43) >= 11'sh0 & $signed(
    inSpriteYPreScaled_43) < 11'sh20 : _GEN_1945; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_44 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_44); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_44_T = $signed(inSpriteXValue_44) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_44_T_4 = inSpriteXValue_44[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_44_T_8 = _inSpriteHorizontal_44_T & $signed(inSpriteXValue_44) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_44_T_5 = {$signed(inSpriteXValue_44), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_44_T_14 = _inSpriteHorizontal_44_T & $signed(inSpriteXValue_44) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1952 = spriteScaleUpHorizontalReg_44 ? $signed({{2{_inSpriteX_44_T_4[10]}},_inSpriteX_44_T_4}) :
    $signed(_inSpriteX_44_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1953 = spriteScaleUpHorizontalReg_44 ? _inSpriteHorizontal_44_T_8 : _inSpriteHorizontal_44_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1954 = ~spriteScaleUpHorizontalReg_44 ? $signed({{1{inSpriteXValue_44[11]}},inSpriteXValue_44}) :
    $signed(_GEN_1952); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_44 = ~spriteScaleUpHorizontalReg_44 ? $signed(inSpriteXValue_44) >= 12'sh0 & $signed(
    inSpriteXValue_44) < 12'sh20 : _GEN_1953; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3439 = {{1{spriteYPositionReg_44[9]}},spriteYPositionReg_44}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_44 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3439); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_44 = inSpriteYValue_44[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_44_T = $signed(inSpriteYPreScaled_44) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_44_T_4 = inSpriteYPreScaled_44[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_44_T_8 = _inSpriteVertical_44_T & $signed(inSpriteYPreScaled_44) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_44_T_5 = {$signed(inSpriteYPreScaled_44), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_44_T_14 = _inSpriteVertical_44_T & $signed(inSpriteYPreScaled_44) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1960 = spriteScaleUpVerticalReg_44 ? $signed({{2{_inSpriteY_44_T_4[9]}},_inSpriteY_44_T_4}) :
    $signed(_inSpriteY_44_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1961 = spriteScaleUpVerticalReg_44 ? _inSpriteVertical_44_T_8 : _inSpriteVertical_44_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1962 = ~spriteScaleUpVerticalReg_44 ? $signed({{1{inSpriteYPreScaled_44[10]}},inSpriteYPreScaled_44})
     : $signed(_GEN_1960); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_44 = ~spriteScaleUpVerticalReg_44 ? $signed(inSpriteYPreScaled_44) >= 11'sh0 & $signed(
    inSpriteYPreScaled_44) < 11'sh20 : _GEN_1961; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_45 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_45); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_45_T = $signed(inSpriteXValue_45) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_45_T_4 = inSpriteXValue_45[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_45_T_8 = _inSpriteHorizontal_45_T & $signed(inSpriteXValue_45) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_45_T_5 = {$signed(inSpriteXValue_45), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_45_T_14 = _inSpriteHorizontal_45_T & $signed(inSpriteXValue_45) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1968 = spriteScaleUpHorizontalReg_45 ? $signed({{2{_inSpriteX_45_T_4[10]}},_inSpriteX_45_T_4}) :
    $signed(_inSpriteX_45_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1969 = spriteScaleUpHorizontalReg_45 ? _inSpriteHorizontal_45_T_8 : _inSpriteHorizontal_45_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1970 = ~spriteScaleUpHorizontalReg_45 ? $signed({{1{inSpriteXValue_45[11]}},inSpriteXValue_45}) :
    $signed(_GEN_1968); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_45 = ~spriteScaleUpHorizontalReg_45 ? $signed(inSpriteXValue_45) >= 12'sh0 & $signed(
    inSpriteXValue_45) < 12'sh20 : _GEN_1969; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3441 = {{1{spriteYPositionReg_45[9]}},spriteYPositionReg_45}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_45 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3441); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_45 = inSpriteYValue_45[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_45_T = $signed(inSpriteYPreScaled_45) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_45_T_4 = inSpriteYPreScaled_45[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_45_T_8 = _inSpriteVertical_45_T & $signed(inSpriteYPreScaled_45) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_45_T_5 = {$signed(inSpriteYPreScaled_45), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_45_T_14 = _inSpriteVertical_45_T & $signed(inSpriteYPreScaled_45) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1976 = spriteScaleUpVerticalReg_45 ? $signed({{2{_inSpriteY_45_T_4[9]}},_inSpriteY_45_T_4}) :
    $signed(_inSpriteY_45_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1977 = spriteScaleUpVerticalReg_45 ? _inSpriteVertical_45_T_8 : _inSpriteVertical_45_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1978 = ~spriteScaleUpVerticalReg_45 ? $signed({{1{inSpriteYPreScaled_45[10]}},inSpriteYPreScaled_45})
     : $signed(_GEN_1976); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_45 = ~spriteScaleUpVerticalReg_45 ? $signed(inSpriteYPreScaled_45) >= 11'sh0 & $signed(
    inSpriteYPreScaled_45) < 11'sh20 : _GEN_1977; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_46 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_46); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_46 = $signed(inSpriteXValue_46) >= 12'sh0 & $signed(inSpriteXValue_46) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1986 = {{1{inSpriteXValue_46[11]}},inSpriteXValue_46}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3443 = {{1{spriteYPositionReg_46[9]}},spriteYPositionReg_46}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_46 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3443); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_46 = inSpriteYValue_46[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_46 = $signed(inSpriteYPreScaled_46) >= 11'sh0 & $signed(inSpriteYPreScaled_46) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1994 = {{1{inSpriteYPreScaled_46[10]}},inSpriteYPreScaled_46}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_47 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_47); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_47 = $signed(inSpriteXValue_47) >= 12'sh0 & $signed(inSpriteXValue_47) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2002 = {{1{inSpriteXValue_47[11]}},inSpriteXValue_47}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3445 = {{1{spriteYPositionReg_47[9]}},spriteYPositionReg_47}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_47 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3445); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_47 = inSpriteYValue_47[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_47 = $signed(inSpriteYPreScaled_47) >= 11'sh0 & $signed(inSpriteYPreScaled_47) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2010 = {{1{inSpriteYPreScaled_47[10]}},inSpriteYPreScaled_47}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_48 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_48); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_48 = $signed(inSpriteXValue_48) >= 12'sh0 & $signed(inSpriteXValue_48) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2018 = {{1{inSpriteXValue_48[11]}},inSpriteXValue_48}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3447 = {{1{spriteYPositionReg_48[9]}},spriteYPositionReg_48}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_48 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3447); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_48 = inSpriteYValue_48[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_48 = $signed(inSpriteYPreScaled_48) >= 11'sh0 & $signed(inSpriteYPreScaled_48) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2026 = {{1{inSpriteYPreScaled_48[10]}},inSpriteYPreScaled_48}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_49 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_49); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_49 = $signed(inSpriteXValue_49) >= 12'sh0 & $signed(inSpriteXValue_49) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2034 = {{1{inSpriteXValue_49[11]}},inSpriteXValue_49}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3449 = {{1{spriteYPositionReg_49[9]}},spriteYPositionReg_49}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_49 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3449); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_49 = inSpriteYValue_49[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_49 = $signed(inSpriteYPreScaled_49) >= 11'sh0 & $signed(inSpriteYPreScaled_49) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2042 = {{1{inSpriteYPreScaled_49[10]}},inSpriteYPreScaled_49}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_50 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_50); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_50 = $signed(inSpriteXValue_50) >= 12'sh0 & $signed(inSpriteXValue_50) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2050 = {{1{inSpriteXValue_50[11]}},inSpriteXValue_50}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3451 = {{1{spriteYPositionReg_50[9]}},spriteYPositionReg_50}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_50 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3451); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_50 = inSpriteYValue_50[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_50 = $signed(inSpriteYPreScaled_50) >= 11'sh0 & $signed(inSpriteYPreScaled_50) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2058 = {{1{inSpriteYPreScaled_50[10]}},inSpriteYPreScaled_50}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_51 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_51); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_51 = $signed(inSpriteXValue_51) >= 12'sh0 & $signed(inSpriteXValue_51) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2066 = {{1{inSpriteXValue_51[11]}},inSpriteXValue_51}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3453 = {{1{spriteYPositionReg_51[9]}},spriteYPositionReg_51}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_51 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3453); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_51 = inSpriteYValue_51[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_51 = $signed(inSpriteYPreScaled_51) >= 11'sh0 & $signed(inSpriteYPreScaled_51) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2074 = {{1{inSpriteYPreScaled_51[10]}},inSpriteYPreScaled_51}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_52 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_52); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_52 = $signed(inSpriteXValue_52) >= 12'sh0 & $signed(inSpriteXValue_52) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2082 = {{1{inSpriteXValue_52[11]}},inSpriteXValue_52}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3455 = {{1{spriteYPositionReg_52[9]}},spriteYPositionReg_52}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_52 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3455); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_52 = inSpriteYValue_52[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_52 = $signed(inSpriteYPreScaled_52) >= 11'sh0 & $signed(inSpriteYPreScaled_52) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2090 = {{1{inSpriteYPreScaled_52[10]}},inSpriteYPreScaled_52}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_53 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_53); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_53 = $signed(inSpriteXValue_53) >= 12'sh0 & $signed(inSpriteXValue_53) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2098 = {{1{inSpriteXValue_53[11]}},inSpriteXValue_53}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3457 = {{1{spriteYPositionReg_53[9]}},spriteYPositionReg_53}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_53 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3457); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_53 = inSpriteYValue_53[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_53 = $signed(inSpriteYPreScaled_53) >= 11'sh0 & $signed(inSpriteYPreScaled_53) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2106 = {{1{inSpriteYPreScaled_53[10]}},inSpriteYPreScaled_53}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_54 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_54); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_54 = $signed(inSpriteXValue_54) >= 12'sh0 & $signed(inSpriteXValue_54) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2114 = {{1{inSpriteXValue_54[11]}},inSpriteXValue_54}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3459 = {{1{spriteYPositionReg_54[9]}},spriteYPositionReg_54}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_54 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3459); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_54 = inSpriteYValue_54[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_54 = $signed(inSpriteYPreScaled_54) >= 11'sh0 & $signed(inSpriteYPreScaled_54) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2122 = {{1{inSpriteYPreScaled_54[10]}},inSpriteYPreScaled_54}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_55 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_55); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_55 = $signed(inSpriteXValue_55) >= 12'sh0 & $signed(inSpriteXValue_55) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2130 = {{1{inSpriteXValue_55[11]}},inSpriteXValue_55}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3461 = {{1{spriteYPositionReg_55[9]}},spriteYPositionReg_55}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_55 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3461); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_55 = inSpriteYValue_55[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_55 = $signed(inSpriteYPreScaled_55) >= 11'sh0 & $signed(inSpriteYPreScaled_55) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2138 = {{1{inSpriteYPreScaled_55[10]}},inSpriteYPreScaled_55}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_56 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_56); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_56 = $signed(inSpriteXValue_56) >= 12'sh0 & $signed(inSpriteXValue_56) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2146 = {{1{inSpriteXValue_56[11]}},inSpriteXValue_56}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3463 = {{1{spriteYPositionReg_56[9]}},spriteYPositionReg_56}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_56 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3463); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_56 = inSpriteYValue_56[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_56 = $signed(inSpriteYPreScaled_56) >= 11'sh0 & $signed(inSpriteYPreScaled_56) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2154 = {{1{inSpriteYPreScaled_56[10]}},inSpriteYPreScaled_56}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_57 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_57); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_57 = $signed(inSpriteXValue_57) >= 12'sh0 & $signed(inSpriteXValue_57) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2162 = {{1{inSpriteXValue_57[11]}},inSpriteXValue_57}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3465 = {{1{spriteYPositionReg_57[9]}},spriteYPositionReg_57}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_57 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3465); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_57 = inSpriteYValue_57[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_57 = $signed(inSpriteYPreScaled_57) >= 11'sh0 & $signed(inSpriteYPreScaled_57) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2170 = {{1{inSpriteYPreScaled_57[10]}},inSpriteYPreScaled_57}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_58 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_58); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_58_T = $signed(inSpriteXValue_58) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_58_T_4 = inSpriteXValue_58[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_58_T_8 = _inSpriteHorizontal_58_T & $signed(inSpriteXValue_58) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_58_T_5 = {$signed(inSpriteXValue_58), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_58_T_14 = _inSpriteHorizontal_58_T & $signed(inSpriteXValue_58) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_2176 = spriteScaleUpHorizontalReg_58 ? $signed({{2{_inSpriteX_58_T_4[10]}},_inSpriteX_58_T_4}) :
    $signed(_inSpriteX_58_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_2177 = spriteScaleUpHorizontalReg_58 ? _inSpriteHorizontal_58_T_8 : _inSpriteHorizontal_58_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_2178 = ~spriteScaleUpHorizontalReg_58 ? $signed({{1{inSpriteXValue_58[11]}},inSpriteXValue_58}) :
    $signed(_GEN_2176); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_58 = ~spriteScaleUpHorizontalReg_58 ? $signed(inSpriteXValue_58) >= 12'sh0 & $signed(
    inSpriteXValue_58) < 12'sh20 : _GEN_2177; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3467 = {{1{spriteYPositionReg_58[9]}},spriteYPositionReg_58}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_58 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3467); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_58 = inSpriteYValue_58[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_58_T = $signed(inSpriteYPreScaled_58) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_58_T_4 = inSpriteYPreScaled_58[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_58_T_8 = _inSpriteVertical_58_T & $signed(inSpriteYPreScaled_58) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_58_T_5 = {$signed(inSpriteYPreScaled_58), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_58_T_14 = _inSpriteVertical_58_T & $signed(inSpriteYPreScaled_58) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_2184 = spriteScaleUpVerticalReg_58 ? $signed({{2{_inSpriteY_58_T_4[9]}},_inSpriteY_58_T_4}) :
    $signed(_inSpriteY_58_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_2185 = spriteScaleUpVerticalReg_58 ? _inSpriteVertical_58_T_8 : _inSpriteVertical_58_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_2186 = ~spriteScaleUpVerticalReg_58 ? $signed({{1{inSpriteYPreScaled_58[10]}},inSpriteYPreScaled_58})
     : $signed(_GEN_2184); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_58 = ~spriteScaleUpVerticalReg_58 ? $signed(inSpriteYPreScaled_58) >= 11'sh0 & $signed(
    inSpriteYPreScaled_58) < 11'sh20 : _GEN_2185; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_59 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_59); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_59_T = $signed(inSpriteXValue_59) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_59_T_4 = inSpriteXValue_59[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_59_T_8 = _inSpriteHorizontal_59_T & $signed(inSpriteXValue_59) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_59_T_5 = {$signed(inSpriteXValue_59), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_59_T_14 = _inSpriteHorizontal_59_T & $signed(inSpriteXValue_59) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_2192 = spriteScaleUpHorizontalReg_59 ? $signed({{2{_inSpriteX_59_T_4[10]}},_inSpriteX_59_T_4}) :
    $signed(_inSpriteX_59_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_2193 = spriteScaleUpHorizontalReg_59 ? _inSpriteHorizontal_59_T_8 : _inSpriteHorizontal_59_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_2194 = ~spriteScaleUpHorizontalReg_59 ? $signed({{1{inSpriteXValue_59[11]}},inSpriteXValue_59}) :
    $signed(_GEN_2192); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_59 = ~spriteScaleUpHorizontalReg_59 ? $signed(inSpriteXValue_59) >= 12'sh0 & $signed(
    inSpriteXValue_59) < 12'sh20 : _GEN_2193; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3469 = {{1{spriteYPositionReg_59[9]}},spriteYPositionReg_59}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_59 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3469); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_59 = inSpriteYValue_59[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_59_T = $signed(inSpriteYPreScaled_59) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_59_T_4 = inSpriteYPreScaled_59[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_59_T_8 = _inSpriteVertical_59_T & $signed(inSpriteYPreScaled_59) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_59_T_5 = {$signed(inSpriteYPreScaled_59), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_59_T_14 = _inSpriteVertical_59_T & $signed(inSpriteYPreScaled_59) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_2200 = spriteScaleUpVerticalReg_59 ? $signed({{2{_inSpriteY_59_T_4[9]}},_inSpriteY_59_T_4}) :
    $signed(_inSpriteY_59_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_2201 = spriteScaleUpVerticalReg_59 ? _inSpriteVertical_59_T_8 : _inSpriteVertical_59_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_2202 = ~spriteScaleUpVerticalReg_59 ? $signed({{1{inSpriteYPreScaled_59[10]}},inSpriteYPreScaled_59})
     : $signed(_GEN_2200); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_59 = ~spriteScaleUpVerticalReg_59 ? $signed(inSpriteYPreScaled_59) >= 11'sh0 & $signed(
    inSpriteYPreScaled_59) < 11'sh20 : _GEN_2201; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_60 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_60); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_60_T = $signed(inSpriteXValue_60) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_60_T_4 = inSpriteXValue_60[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_60_T_8 = _inSpriteHorizontal_60_T & $signed(inSpriteXValue_60) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_60_T_5 = {$signed(inSpriteXValue_60), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_60_T_14 = _inSpriteHorizontal_60_T & $signed(inSpriteXValue_60) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_2208 = spriteScaleUpHorizontalReg_60 ? $signed({{2{_inSpriteX_60_T_4[10]}},_inSpriteX_60_T_4}) :
    $signed(_inSpriteX_60_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_2209 = spriteScaleUpHorizontalReg_60 ? _inSpriteHorizontal_60_T_8 : _inSpriteHorizontal_60_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_2210 = ~spriteScaleUpHorizontalReg_60 ? $signed({{1{inSpriteXValue_60[11]}},inSpriteXValue_60}) :
    $signed(_GEN_2208); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_60 = ~spriteScaleUpHorizontalReg_60 ? $signed(inSpriteXValue_60) >= 12'sh0 & $signed(
    inSpriteXValue_60) < 12'sh20 : _GEN_2209; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_3471 = {{1{spriteYPositionReg_60[9]}},spriteYPositionReg_60}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_60 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3471); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_60 = inSpriteYValue_60[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_60_T = $signed(inSpriteYPreScaled_60) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_60_T_4 = inSpriteYPreScaled_60[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_60_T_8 = _inSpriteVertical_60_T & $signed(inSpriteYPreScaled_60) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_60_T_5 = {$signed(inSpriteYPreScaled_60), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_60_T_14 = _inSpriteVertical_60_T & $signed(inSpriteYPreScaled_60) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_2216 = spriteScaleUpVerticalReg_60 ? $signed({{2{_inSpriteY_60_T_4[9]}},_inSpriteY_60_T_4}) :
    $signed(_inSpriteY_60_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_2217 = spriteScaleUpVerticalReg_60 ? _inSpriteVertical_60_T_8 : _inSpriteVertical_60_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_2218 = ~spriteScaleUpVerticalReg_60 ? $signed({{1{inSpriteYPreScaled_60[10]}},inSpriteYPreScaled_60})
     : $signed(_GEN_2216); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_60 = ~spriteScaleUpVerticalReg_60 ? $signed(inSpriteYPreScaled_60) >= 11'sh0 & $signed(
    inSpriteYPreScaled_60) < 11'sh20 : _GEN_2217; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_61 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_61); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_61 = $signed(inSpriteXValue_61) >= 12'sh0 & $signed(inSpriteXValue_61) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2226 = {{1{inSpriteXValue_61[11]}},inSpriteXValue_61}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3473 = {{1{spriteYPositionReg_61[9]}},spriteYPositionReg_61}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_61 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3473); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_61 = inSpriteYValue_61[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_61 = $signed(inSpriteYPreScaled_61) >= 11'sh0 & $signed(inSpriteYPreScaled_61) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2234 = {{1{inSpriteYPreScaled_61[10]}},inSpriteYPreScaled_61}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_62 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_62); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_62 = $signed(inSpriteXValue_62) >= 12'sh0 & $signed(inSpriteXValue_62) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2242 = {{1{inSpriteXValue_62[11]}},inSpriteXValue_62}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3475 = {{1{spriteYPositionReg_62[9]}},spriteYPositionReg_62}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_62 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3475); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_62 = inSpriteYValue_62[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_62 = $signed(inSpriteYPreScaled_62) >= 11'sh0 & $signed(inSpriteYPreScaled_62) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2250 = {{1{inSpriteYPreScaled_62[10]}},inSpriteYPreScaled_62}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_63 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_63); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_63 = $signed(inSpriteXValue_63) >= 12'sh0 & $signed(inSpriteXValue_63) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_2258 = {{1{inSpriteXValue_63[11]}},inSpriteXValue_63}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_3477 = {{1{spriteYPositionReg_63[9]}},spriteYPositionReg_63}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_63 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_3477); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_63 = inSpriteYValue_63[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_63 = $signed(inSpriteYPreScaled_63) >= 11'sh0 & $signed(inSpriteYPreScaled_63) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_2266 = {{1{inSpriteYPreScaled_63[10]}},inSpriteYPreScaled_63}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteX_0 = _GEN_1250[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_0 = _GEN_1258[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_0_io_address_T_2 = 6'h20 * inSpriteY_0[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3545 = {{6'd0}, inSpriteX_0[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_0_io_address_T_4 = _GEN_3545 + _spriteMemories_0_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_3 = _GEN_1298[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_3 = _GEN_1306[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_3_io_address_T_2 = 6'h20 * inSpriteY_3[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3554 = {{6'd0}, inSpriteX_3[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_3_io_address_T_4 = _GEN_3554 + _spriteMemories_3_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_7 = _GEN_1362[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_7 = _GEN_1370[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_7_io_address_T_2 = 6'h20 * inSpriteY_7[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3566 = {{6'd0}, inSpriteX_7[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_7_io_address_T_4 = _GEN_3566 + _spriteMemories_7_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_8 = _GEN_1378[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_8 = _GEN_1386[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_8_io_address_T_2 = 6'h20 * inSpriteY_8[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3569 = {{6'd0}, inSpriteX_8[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_8_io_address_T_4 = _GEN_3569 + _spriteMemories_8_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_9 = _GEN_1394[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_9 = _GEN_1402[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_9_io_address_T_2 = 6'h20 * inSpriteY_9[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3572 = {{6'd0}, inSpriteX_9[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_9_io_address_T_4 = _GEN_3572 + _spriteMemories_9_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_10 = _GEN_1410[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_10 = _GEN_1418[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_10_io_address_T_2 = 6'h20 * inSpriteY_10[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3575 = {{6'd0}, inSpriteX_10[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_10_io_address_T_4 = _GEN_3575 + _spriteMemories_10_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_11 = _GEN_1426[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_11 = _GEN_1434[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_11_io_address_T_2 = 6'h20 * inSpriteY_11[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3578 = {{6'd0}, inSpriteX_11[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_11_io_address_T_4 = _GEN_3578 + _spriteMemories_11_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_12 = _GEN_1442[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_12 = _GEN_1450[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_12_io_address_T_2 = 6'h20 * inSpriteY_12[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3581 = {{6'd0}, inSpriteX_12[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_12_io_address_T_4 = _GEN_3581 + _spriteMemories_12_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_13 = _GEN_1458[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_13 = _GEN_1466[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_13_io_address_T_2 = 6'h20 * inSpriteY_13[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3584 = {{6'd0}, inSpriteX_13[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_13_io_address_T_4 = _GEN_3584 + _spriteMemories_13_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_14 = _GEN_1474[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_14 = _GEN_1482[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_14_io_address_T_2 = 6'h20 * inSpriteY_14[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3587 = {{6'd0}, inSpriteX_14[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_14_io_address_T_4 = _GEN_3587 + _spriteMemories_14_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_16 = _GEN_1506[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_16 = _GEN_1514[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_16_io_address_T_2 = 6'h20 * inSpriteY_16[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3593 = {{6'd0}, inSpriteX_16[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_16_io_address_T_4 = _GEN_3593 + _spriteMemories_16_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_17 = _GEN_1522[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_17 = _GEN_1530[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_17_io_address_T_2 = 6'h20 * inSpriteY_17[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3596 = {{6'd0}, inSpriteX_17[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_17_io_address_T_4 = _GEN_3596 + _spriteMemories_17_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_18 = _GEN_1538[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_18 = _GEN_1546[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_18_io_address_T_2 = 6'h20 * inSpriteY_18[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3599 = {{6'd0}, inSpriteX_18[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_18_io_address_T_4 = _GEN_3599 + _spriteMemories_18_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_19 = _GEN_1554[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_19 = _GEN_1562[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_19_io_address_T_2 = 6'h20 * inSpriteY_19[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3602 = {{6'd0}, inSpriteX_19[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_19_io_address_T_4 = _GEN_3602 + _spriteMemories_19_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_20 = _GEN_1570[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_20 = _GEN_1578[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_20_io_address_T_2 = 6'h20 * inSpriteY_20[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3605 = {{6'd0}, inSpriteX_20[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_20_io_address_T_4 = _GEN_3605 + _spriteMemories_20_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_21 = _GEN_1586[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_21 = _GEN_1594[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_21_io_address_T_2 = 6'h20 * inSpriteY_21[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3608 = {{6'd0}, inSpriteX_21[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_21_io_address_T_4 = _GEN_3608 + _spriteMemories_21_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_22 = _GEN_1602[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_22 = _GEN_1610[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_22_io_address_T_2 = 6'h20 * inSpriteY_22[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3611 = {{6'd0}, inSpriteX_22[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_22_io_address_T_4 = _GEN_3611 + _spriteMemories_22_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_23 = _GEN_1618[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_23 = _GEN_1626[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_23_io_address_T_2 = 6'h20 * inSpriteY_23[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3614 = {{6'd0}, inSpriteX_23[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_23_io_address_T_4 = _GEN_3614 + _spriteMemories_23_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_24 = _GEN_1634[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_24 = _GEN_1642[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_24_io_address_T_2 = 6'h20 * inSpriteY_24[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3617 = {{6'd0}, inSpriteX_24[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_24_io_address_T_4 = _GEN_3617 + _spriteMemories_24_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_25 = _GEN_1650[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_25 = _GEN_1658[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_25_io_address_T_2 = 6'h20 * inSpriteY_25[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3620 = {{6'd0}, inSpriteX_25[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_25_io_address_T_4 = _GEN_3620 + _spriteMemories_25_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_26 = _GEN_1666[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_26 = _GEN_1674[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_26_io_address_T_2 = 6'h20 * inSpriteY_26[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3623 = {{6'd0}, inSpriteX_26[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_26_io_address_T_4 = _GEN_3623 + _spriteMemories_26_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_27 = _GEN_1682[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_27 = _GEN_1690[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_27_io_address_T_2 = 6'h20 * inSpriteY_27[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3626 = {{6'd0}, inSpriteX_27[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_27_io_address_T_4 = _GEN_3626 + _spriteMemories_27_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_28 = _GEN_1698[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_28 = _GEN_1706[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_28_io_address_T_2 = 6'h20 * inSpriteY_28[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3629 = {{6'd0}, inSpriteX_28[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_28_io_address_T_4 = _GEN_3629 + _spriteMemories_28_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_29 = _GEN_1714[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_29 = _GEN_1722[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_29_io_address_T_2 = 6'h20 * inSpriteY_29[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3632 = {{6'd0}, inSpriteX_29[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_29_io_address_T_4 = _GEN_3632 + _spriteMemories_29_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_30 = _GEN_1730[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_30 = _GEN_1738[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_30_io_address_T_2 = 6'h20 * inSpriteY_30[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3635 = {{6'd0}, inSpriteX_30[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_30_io_address_T_4 = _GEN_3635 + _spriteMemories_30_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_31 = _GEN_1746[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_31 = _GEN_1754[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_31_io_address_T_2 = 6'h20 * inSpriteY_31[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3638 = {{6'd0}, inSpriteX_31[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_31_io_address_T_4 = _GEN_3638 + _spriteMemories_31_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_32 = _GEN_1762[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_32 = _GEN_1770[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_32_io_address_T_2 = 6'h20 * inSpriteY_32[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3641 = {{6'd0}, inSpriteX_32[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_32_io_address_T_4 = _GEN_3641 + _spriteMemories_32_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_33 = _GEN_1778[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_33 = _GEN_1786[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_33_io_address_T_2 = 6'h20 * inSpriteY_33[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3644 = {{6'd0}, inSpriteX_33[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_33_io_address_T_4 = _GEN_3644 + _spriteMemories_33_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_34 = _GEN_1794[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_34 = _GEN_1802[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_34_io_address_T_2 = 6'h20 * inSpriteY_34[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3647 = {{6'd0}, inSpriteX_34[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_34_io_address_T_4 = _GEN_3647 + _spriteMemories_34_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_35 = _GEN_1810[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_35 = _GEN_1818[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_35_io_address_T_2 = 6'h20 * inSpriteY_35[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3650 = {{6'd0}, inSpriteX_35[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_35_io_address_T_4 = _GEN_3650 + _spriteMemories_35_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_36 = _GEN_1826[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_36 = _GEN_1834[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_36_io_address_T_2 = 6'h20 * inSpriteY_36[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3653 = {{6'd0}, inSpriteX_36[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_36_io_address_T_4 = _GEN_3653 + _spriteMemories_36_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_37 = _GEN_1842[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_37 = _GEN_1850[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_37_io_address_T_2 = 6'h20 * inSpriteY_37[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3656 = {{6'd0}, inSpriteX_37[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_37_io_address_T_4 = _GEN_3656 + _spriteMemories_37_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_38 = _GEN_1858[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_38 = _GEN_1866[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_38_io_address_T_2 = 6'h20 * inSpriteY_38[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3659 = {{6'd0}, inSpriteX_38[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_38_io_address_T_4 = _GEN_3659 + _spriteMemories_38_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_39 = _GEN_1874[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_39 = _GEN_1882[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_39_io_address_T_2 = 6'h20 * inSpriteY_39[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3662 = {{6'd0}, inSpriteX_39[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_39_io_address_T_4 = _GEN_3662 + _spriteMemories_39_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_40 = _GEN_1890[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_40 = _GEN_1898[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_40_io_address_T_2 = 6'h20 * inSpriteY_40[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3665 = {{6'd0}, inSpriteX_40[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_40_io_address_T_4 = _GEN_3665 + _spriteMemories_40_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_41 = _GEN_1906[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_41 = _GEN_1914[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_41_io_address_T_2 = 6'h20 * inSpriteY_41[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3668 = {{6'd0}, inSpriteX_41[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_41_io_address_T_4 = _GEN_3668 + _spriteMemories_41_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_42 = _GEN_1922[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_42 = _GEN_1930[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_42_io_address_T_2 = 6'h20 * inSpriteY_42[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3671 = {{6'd0}, inSpriteX_42[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_42_io_address_T_4 = _GEN_3671 + _spriteMemories_42_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_43 = _GEN_1938[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_43 = _GEN_1946[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_43_io_address_T_2 = 6'h20 * inSpriteY_43[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3674 = {{6'd0}, inSpriteX_43[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_43_io_address_T_4 = _GEN_3674 + _spriteMemories_43_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_44 = _GEN_1954[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_44 = _GEN_1962[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_44_io_address_T_2 = 6'h20 * inSpriteY_44[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3677 = {{6'd0}, inSpriteX_44[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_44_io_address_T_4 = _GEN_3677 + _spriteMemories_44_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_45 = _GEN_1970[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_45 = _GEN_1978[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_45_io_address_T_2 = 6'h20 * inSpriteY_45[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3680 = {{6'd0}, inSpriteX_45[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_45_io_address_T_4 = _GEN_3680 + _spriteMemories_45_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_46 = _GEN_1986[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_46 = _GEN_1994[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_46_io_address_T_2 = 6'h20 * inSpriteY_46[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3683 = {{6'd0}, inSpriteX_46[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_46_io_address_T_4 = _GEN_3683 + _spriteMemories_46_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_47 = _GEN_2002[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_47 = _GEN_2010[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_47_io_address_T_2 = 6'h20 * inSpriteY_47[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3686 = {{6'd0}, inSpriteX_47[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_47_io_address_T_4 = _GEN_3686 + _spriteMemories_47_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_48 = _GEN_2018[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_48 = _GEN_2026[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_48_io_address_T_2 = 6'h20 * inSpriteY_48[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3689 = {{6'd0}, inSpriteX_48[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_48_io_address_T_4 = _GEN_3689 + _spriteMemories_48_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_49 = _GEN_2034[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_49 = _GEN_2042[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_49_io_address_T_2 = 6'h20 * inSpriteY_49[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3692 = {{6'd0}, inSpriteX_49[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_49_io_address_T_4 = _GEN_3692 + _spriteMemories_49_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_50 = _GEN_2050[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_50 = _GEN_2058[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_50_io_address_T_2 = 6'h20 * inSpriteY_50[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3695 = {{6'd0}, inSpriteX_50[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_50_io_address_T_4 = _GEN_3695 + _spriteMemories_50_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_51 = _GEN_2066[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_51 = _GEN_2074[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_51_io_address_T_2 = 6'h20 * inSpriteY_51[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3698 = {{6'd0}, inSpriteX_51[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_51_io_address_T_4 = _GEN_3698 + _spriteMemories_51_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_52 = _GEN_2082[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_52 = _GEN_2090[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_52_io_address_T_2 = 6'h20 * inSpriteY_52[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3701 = {{6'd0}, inSpriteX_52[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_52_io_address_T_4 = _GEN_3701 + _spriteMemories_52_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_53 = _GEN_2098[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_53 = _GEN_2106[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_53_io_address_T_2 = 6'h20 * inSpriteY_53[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3704 = {{6'd0}, inSpriteX_53[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_53_io_address_T_4 = _GEN_3704 + _spriteMemories_53_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_54 = _GEN_2114[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_54 = _GEN_2122[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_54_io_address_T_2 = 6'h20 * inSpriteY_54[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3707 = {{6'd0}, inSpriteX_54[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_54_io_address_T_4 = _GEN_3707 + _spriteMemories_54_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_55 = _GEN_2130[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_55 = _GEN_2138[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_55_io_address_T_2 = 6'h20 * inSpriteY_55[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3710 = {{6'd0}, inSpriteX_55[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_55_io_address_T_4 = _GEN_3710 + _spriteMemories_55_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_56 = _GEN_2146[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_56 = _GEN_2154[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_56_io_address_T_2 = 6'h20 * inSpriteY_56[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3713 = {{6'd0}, inSpriteX_56[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_56_io_address_T_4 = _GEN_3713 + _spriteMemories_56_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_57 = _GEN_2162[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_57 = _GEN_2170[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_57_io_address_T_2 = 6'h20 * inSpriteY_57[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3716 = {{6'd0}, inSpriteX_57[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_57_io_address_T_4 = _GEN_3716 + _spriteMemories_57_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_58 = _GEN_2178[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_58 = _GEN_2186[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_58_io_address_T_2 = 6'h20 * inSpriteY_58[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3719 = {{6'd0}, inSpriteX_58[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_58_io_address_T_4 = _GEN_3719 + _spriteMemories_58_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_59 = _GEN_2194[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_59 = _GEN_2202[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_59_io_address_T_2 = 6'h20 * inSpriteY_59[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3722 = {{6'd0}, inSpriteX_59[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_59_io_address_T_4 = _GEN_3722 + _spriteMemories_59_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_60 = _GEN_2210[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_60 = _GEN_2218[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_60_io_address_T_2 = 6'h20 * inSpriteY_60[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3725 = {{6'd0}, inSpriteX_60[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_60_io_address_T_4 = _GEN_3725 + _spriteMemories_60_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_61 = _GEN_2226[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_61 = _GEN_2234[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_61_io_address_T_2 = 6'h20 * inSpriteY_61[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3728 = {{6'd0}, inSpriteX_61[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_61_io_address_T_4 = _GEN_3728 + _spriteMemories_61_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_62 = _GEN_2242[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_62 = _GEN_2250[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_62_io_address_T_2 = 6'h20 * inSpriteY_62[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3731 = {{6'd0}, inSpriteX_62[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_62_io_address_T_4 = _GEN_3731 + _spriteMemories_62_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_63 = _GEN_2258[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_63 = _GEN_2266[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_63_io_address_T_2 = 6'h20 * inSpriteY_63[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_3734 = {{6'd0}, inSpriteX_63[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_63_io_address_T_4 = _GEN_3734 + _spriteMemories_63_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_64_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_64_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_64_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_64_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_64_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_64_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_65_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_65_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_65_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_65_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_65_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_65_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_66_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_66_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_66_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_66_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_66_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_66_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_67_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_67_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_67_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_67_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_67_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_67_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_68_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_68_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_68_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_68_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_68_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_68_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_69_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_69_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_69_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_69_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_69_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_69_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_70_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_70_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_70_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_70_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_70_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_70_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_71_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_71_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_71_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_71_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_71_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_71_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_72_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_72_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_72_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_72_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_72_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_72_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_73_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_73_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_73_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_73_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_73_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_73_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_74_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_74_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_74_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_74_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_74_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_74_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_75_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_75_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_75_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_75_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_75_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_75_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_76_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_76_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_76_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_76_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_76_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_76_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_77_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_77_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_77_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_77_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_77_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_77_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_78_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_78_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_78_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_78_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_78_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_78_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_79_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_79_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_79_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_79_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_79_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_79_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_80_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_80_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_80_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_80_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_80_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_80_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_81_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_81_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_81_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_81_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_81_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_81_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_82_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_82_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_82_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_82_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_82_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_82_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_83_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_83_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_83_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_83_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_83_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_83_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_84_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_84_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_84_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_84_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_84_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_84_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_85_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_85_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_85_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_85_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_85_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_85_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_86_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_86_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_86_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_86_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_86_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_86_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_87_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_87_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_87_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_87_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_87_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_87_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_88_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_88_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_88_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_88_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_88_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_88_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_89_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_89_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_89_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_89_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_89_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_89_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_90_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_90_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_90_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_90_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_90_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_90_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_91_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_91_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_91_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_91_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_91_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_91_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_92_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_92_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_92_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_92_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_92_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_92_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_93_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_93_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_93_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_93_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_93_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_93_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_94_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_94_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_94_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_94_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_94_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_94_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_95_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_95_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_95_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_95_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_95_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_95_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_96_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_96_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_96_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_96_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_96_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_96_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_97_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_97_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_97_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_97_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_97_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_97_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_98_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_98_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_98_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_98_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_98_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_98_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_99_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_99_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_99_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_99_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_99_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_99_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_100_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_100_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_100_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_100_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_100_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_100_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_101_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_101_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_101_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_101_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_101_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_101_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_102_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_102_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_102_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_102_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_102_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_102_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_103_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_103_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_103_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_103_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_103_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_103_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_104_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_104_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_104_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_104_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_104_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_104_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_105_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_105_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_105_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_105_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_105_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_105_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_106_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_106_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_106_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_106_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_106_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_106_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_107_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_107_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_107_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_107_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_107_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_107_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_108_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_108_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_108_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_108_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_108_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_108_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_109_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_109_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_109_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_109_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_109_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_109_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_110_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_110_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_110_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_110_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_110_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_110_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_111_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_111_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_111_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_111_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_111_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_111_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_112_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_112_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_112_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_112_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_112_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_112_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_113_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_113_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_113_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_113_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_113_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_113_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_114_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_114_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_114_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_114_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_114_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_114_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_115_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_115_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_115_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_115_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_115_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_115_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_116_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_116_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_116_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_116_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_116_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_116_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_117_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_117_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_117_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_117_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_117_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_117_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_118_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_118_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_118_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_118_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_118_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_118_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_119_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_119_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_119_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_119_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_119_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_119_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_120_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_120_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_120_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_120_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_120_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_120_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_121_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_121_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_121_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_121_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_121_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_121_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_122_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_122_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_122_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_122_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_122_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_122_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_123_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_123_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_123_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_123_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_123_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_123_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_124_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_124_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_124_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_124_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_124_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_124_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_125_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_125_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_125_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_125_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_125_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_125_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_126_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_126_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_126_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_126_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_126_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_126_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_127_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_127_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_127_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_127_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_127_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_127_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] pixelColorSprite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 339:33]
  reg  pixelColorSpriteValid; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 340:38]
  wire [5:0] pixelColorInDisplay = pixelColorSpriteValid ? pixelColorSprite : pixelColorBack; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 344:32]
  reg  pixelColourVGA_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  pixelColourVGA_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  pixelColourVGA_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  wire [5:0] pixelColourVGA = pixelColourVGA_pipeReg_0 ? pixelColorInDisplay : 6'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 345:27]
  reg [3:0] io_vgaRed_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 349:23]
  reg [3:0] io_vgaGreen_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 350:25]
  reg [3:0] io_vgaBlue_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 351:24]
  Memory backTileMemories_0 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_0_clock),
    .io_address(backTileMemories_0_io_address),
    .io_dataRead(backTileMemories_0_io_dataRead)
  );
  Memory_1 backTileMemories_1 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_1_clock),
    .io_address(backTileMemories_1_io_address),
    .io_dataRead(backTileMemories_1_io_dataRead)
  );
  Memory_2 backTileMemories_2 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_2_clock),
    .io_address(backTileMemories_2_io_address),
    .io_dataRead(backTileMemories_2_io_dataRead)
  );
  Memory_3 backTileMemories_3 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_3_clock),
    .io_address(backTileMemories_3_io_address),
    .io_dataRead(backTileMemories_3_io_dataRead)
  );
  Memory_4 backTileMemories_4 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_4_clock),
    .io_address(backTileMemories_4_io_address),
    .io_dataRead(backTileMemories_4_io_dataRead)
  );
  Memory_5 backTileMemories_5 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_5_clock),
    .io_address(backTileMemories_5_io_address),
    .io_dataRead(backTileMemories_5_io_dataRead)
  );
  Memory_6 backTileMemories_6 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_6_clock),
    .io_address(backTileMemories_6_io_address),
    .io_dataRead(backTileMemories_6_io_dataRead)
  );
  Memory_7 backTileMemories_7 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_7_clock),
    .io_address(backTileMemories_7_io_address),
    .io_dataRead(backTileMemories_7_io_dataRead)
  );
  Memory_8 backTileMemories_8 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_8_clock),
    .io_address(backTileMemories_8_io_address),
    .io_dataRead(backTileMemories_8_io_dataRead)
  );
  Memory_9 backTileMemories_9 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_9_clock),
    .io_address(backTileMemories_9_io_address),
    .io_dataRead(backTileMemories_9_io_dataRead)
  );
  Memory_10 backTileMemories_10 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_10_clock),
    .io_address(backTileMemories_10_io_address),
    .io_dataRead(backTileMemories_10_io_dataRead)
  );
  Memory_11 backTileMemories_11 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_11_clock),
    .io_address(backTileMemories_11_io_address),
    .io_dataRead(backTileMemories_11_io_dataRead)
  );
  Memory_12 backTileMemories_12 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_12_clock),
    .io_address(backTileMemories_12_io_address),
    .io_dataRead(backTileMemories_12_io_dataRead)
  );
  Memory_13 backTileMemories_13 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_13_clock),
    .io_address(backTileMemories_13_io_address),
    .io_dataRead(backTileMemories_13_io_dataRead)
  );
  Memory_14 backTileMemories_14 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_14_clock),
    .io_address(backTileMemories_14_io_address),
    .io_dataRead(backTileMemories_14_io_dataRead)
  );
  Memory_15 backTileMemories_15 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_15_clock),
    .io_address(backTileMemories_15_io_address),
    .io_dataRead(backTileMemories_15_io_dataRead)
  );
  Memory_16 backTileMemories_16 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_16_clock),
    .io_address(backTileMemories_16_io_address),
    .io_dataRead(backTileMemories_16_io_dataRead)
  );
  Memory_17 backTileMemories_17 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_17_clock),
    .io_address(backTileMemories_17_io_address),
    .io_dataRead(backTileMemories_17_io_dataRead)
  );
  Memory_18 backTileMemories_18 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_18_clock),
    .io_address(backTileMemories_18_io_address),
    .io_dataRead(backTileMemories_18_io_dataRead)
  );
  Memory_19 backTileMemories_19 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_19_clock),
    .io_address(backTileMemories_19_io_address),
    .io_dataRead(backTileMemories_19_io_dataRead)
  );
  Memory_20 backTileMemories_20 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_20_clock),
    .io_address(backTileMemories_20_io_address),
    .io_dataRead(backTileMemories_20_io_dataRead)
  );
  Memory_21 backTileMemories_21 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_21_clock),
    .io_address(backTileMemories_21_io_address),
    .io_dataRead(backTileMemories_21_io_dataRead)
  );
  Memory_22 backTileMemories_22 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_22_clock),
    .io_address(backTileMemories_22_io_address),
    .io_dataRead(backTileMemories_22_io_dataRead)
  );
  Memory_23 backTileMemories_23 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_23_clock),
    .io_address(backTileMemories_23_io_address),
    .io_dataRead(backTileMemories_23_io_dataRead)
  );
  Memory_24 backTileMemories_24 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_24_clock),
    .io_address(backTileMemories_24_io_address),
    .io_dataRead(backTileMemories_24_io_dataRead)
  );
  Memory_25 backTileMemories_25 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_25_clock),
    .io_address(backTileMemories_25_io_address),
    .io_dataRead(backTileMemories_25_io_dataRead)
  );
  Memory_26 backTileMemories_26 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_26_clock),
    .io_address(backTileMemories_26_io_address),
    .io_dataRead(backTileMemories_26_io_dataRead)
  );
  Memory_27 backTileMemories_27 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_27_clock),
    .io_address(backTileMemories_27_io_address),
    .io_dataRead(backTileMemories_27_io_dataRead)
  );
  Memory_28 backTileMemories_28 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_28_clock),
    .io_address(backTileMemories_28_io_address),
    .io_dataRead(backTileMemories_28_io_dataRead)
  );
  Memory_29 backTileMemories_29 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_29_clock),
    .io_address(backTileMemories_29_io_address),
    .io_dataRead(backTileMemories_29_io_dataRead)
  );
  Memory_30 backTileMemories_30 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_30_clock),
    .io_address(backTileMemories_30_io_address),
    .io_dataRead(backTileMemories_30_io_dataRead)
  );
  Memory_31 backTileMemories_31 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_31_clock),
    .io_address(backTileMemories_31_io_address),
    .io_dataRead(backTileMemories_31_io_dataRead)
  );
  Memory_32 backTileMemories_32 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_32_clock),
    .io_address(backTileMemories_32_io_address),
    .io_dataRead(backTileMemories_32_io_dataRead)
  );
  Memory_33 backTileMemories_33 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_33_clock),
    .io_address(backTileMemories_33_io_address),
    .io_dataRead(backTileMemories_33_io_dataRead)
  );
  Memory_34 backTileMemories_34 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_34_clock),
    .io_address(backTileMemories_34_io_address),
    .io_dataRead(backTileMemories_34_io_dataRead)
  );
  Memory_35 backTileMemories_35 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_35_clock),
    .io_address(backTileMemories_35_io_address),
    .io_dataRead(backTileMemories_35_io_dataRead)
  );
  Memory_36 backTileMemories_36 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_36_clock),
    .io_address(backTileMemories_36_io_address),
    .io_dataRead(backTileMemories_36_io_dataRead)
  );
  Memory_37 backTileMemories_37 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_37_clock),
    .io_address(backTileMemories_37_io_address),
    .io_dataRead(backTileMemories_37_io_dataRead)
  );
  Memory_38 backTileMemories_38 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_38_clock),
    .io_address(backTileMemories_38_io_address),
    .io_dataRead(backTileMemories_38_io_dataRead)
  );
  Memory_39 backTileMemories_39 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_39_clock),
    .io_address(backTileMemories_39_io_address),
    .io_dataRead(backTileMemories_39_io_dataRead)
  );
  Memory_40 backTileMemories_40 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_40_clock),
    .io_address(backTileMemories_40_io_address),
    .io_dataRead(backTileMemories_40_io_dataRead)
  );
  Memory_41 backTileMemories_41 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_41_clock),
    .io_address(backTileMemories_41_io_address),
    .io_dataRead(backTileMemories_41_io_dataRead)
  );
  Memory_42 backTileMemories_42 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_42_clock),
    .io_address(backTileMemories_42_io_address),
    .io_dataRead(backTileMemories_42_io_dataRead)
  );
  Memory_43 backTileMemories_43 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_43_clock),
    .io_address(backTileMemories_43_io_address),
    .io_dataRead(backTileMemories_43_io_dataRead)
  );
  Memory_44 backTileMemories_44 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_44_clock),
    .io_address(backTileMemories_44_io_address),
    .io_dataRead(backTileMemories_44_io_dataRead)
  );
  Memory_45 backTileMemories_45 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_45_clock),
    .io_address(backTileMemories_45_io_address),
    .io_dataRead(backTileMemories_45_io_dataRead)
  );
  Memory_46 backTileMemories_46 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_46_clock),
    .io_address(backTileMemories_46_io_address),
    .io_dataRead(backTileMemories_46_io_dataRead)
  );
  Memory_47 backTileMemories_47 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_47_clock),
    .io_address(backTileMemories_47_io_address),
    .io_dataRead(backTileMemories_47_io_dataRead)
  );
  Memory_48 backTileMemories_48 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_48_clock),
    .io_address(backTileMemories_48_io_address),
    .io_dataRead(backTileMemories_48_io_dataRead)
  );
  Memory_49 backTileMemories_49 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_49_clock),
    .io_address(backTileMemories_49_io_address),
    .io_dataRead(backTileMemories_49_io_dataRead)
  );
  Memory_50 backTileMemories_50 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_50_clock),
    .io_address(backTileMemories_50_io_address),
    .io_dataRead(backTileMemories_50_io_dataRead)
  );
  Memory_51 backTileMemories_51 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_51_clock),
    .io_address(backTileMemories_51_io_address),
    .io_dataRead(backTileMemories_51_io_dataRead)
  );
  Memory_52 backTileMemories_52 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_52_clock),
    .io_address(backTileMemories_52_io_address),
    .io_dataRead(backTileMemories_52_io_dataRead)
  );
  Memory_53 backTileMemories_53 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_53_clock),
    .io_address(backTileMemories_53_io_address),
    .io_dataRead(backTileMemories_53_io_dataRead)
  );
  Memory_54 backTileMemories_54 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_54_clock),
    .io_address(backTileMemories_54_io_address),
    .io_dataRead(backTileMemories_54_io_dataRead)
  );
  Memory_55 backTileMemories_55 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_55_clock),
    .io_address(backTileMemories_55_io_address),
    .io_dataRead(backTileMemories_55_io_dataRead)
  );
  Memory_56 backTileMemories_56 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_56_clock),
    .io_address(backTileMemories_56_io_address),
    .io_dataRead(backTileMemories_56_io_dataRead)
  );
  Memory_57 backTileMemories_57 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_57_clock),
    .io_address(backTileMemories_57_io_address),
    .io_dataRead(backTileMemories_57_io_dataRead)
  );
  Memory_58 backTileMemories_58 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_58_clock),
    .io_address(backTileMemories_58_io_address),
    .io_dataRead(backTileMemories_58_io_dataRead)
  );
  Memory_59 backTileMemories_59 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_59_clock),
    .io_address(backTileMemories_59_io_address),
    .io_dataRead(backTileMemories_59_io_dataRead)
  );
  Memory_60 backTileMemories_60 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_60_clock),
    .io_address(backTileMemories_60_io_address),
    .io_dataRead(backTileMemories_60_io_dataRead)
  );
  Memory_61 backTileMemories_61 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_61_clock),
    .io_address(backTileMemories_61_io_address),
    .io_dataRead(backTileMemories_61_io_dataRead)
  );
  Memory_62 backTileMemories_62 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_62_clock),
    .io_address(backTileMemories_62_io_address),
    .io_dataRead(backTileMemories_62_io_dataRead)
  );
  Memory_63 backTileMemories_63 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_63_clock),
    .io_address(backTileMemories_63_io_address),
    .io_dataRead(backTileMemories_63_io_dataRead)
  );
  Memory_64 backBufferMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
    .clock(backBufferMemory_clock),
    .io_address(backBufferMemory_io_address),
    .io_dataRead(backBufferMemory_io_dataRead),
    .io_writeEnable(backBufferMemory_io_writeEnable),
    .io_dataWrite(backBufferMemory_io_dataWrite)
  );
  Memory_64 backBufferShadowMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
    .clock(backBufferShadowMemory_clock),
    .io_address(backBufferShadowMemory_io_address),
    .io_dataRead(backBufferShadowMemory_io_dataRead),
    .io_writeEnable(backBufferShadowMemory_io_writeEnable),
    .io_dataWrite(backBufferShadowMemory_io_dataWrite)
  );
  Memory_66 backBufferRestoreMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
    .clock(backBufferRestoreMemory_clock),
    .io_address(backBufferRestoreMemory_io_address),
    .io_dataRead(backBufferRestoreMemory_io_dataRead)
  );
  Memory_67 spriteMemories_0 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_0_clock),
    .io_address(spriteMemories_0_io_address),
    .io_dataRead(spriteMemories_0_io_dataRead)
  );
  Memory_68 spriteMemories_1 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_1_clock),
    .io_address(spriteMemories_1_io_address),
    .io_dataRead(spriteMemories_1_io_dataRead)
  );
  Memory_69 spriteMemories_2 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_2_clock),
    .io_address(spriteMemories_2_io_address),
    .io_dataRead(spriteMemories_2_io_dataRead)
  );
  Memory_70 spriteMemories_3 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_3_clock),
    .io_address(spriteMemories_3_io_address),
    .io_dataRead(spriteMemories_3_io_dataRead)
  );
  Memory_71 spriteMemories_4 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_4_clock),
    .io_address(spriteMemories_4_io_address),
    .io_dataRead(spriteMemories_4_io_dataRead)
  );
  Memory_72 spriteMemories_5 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_5_clock),
    .io_address(spriteMemories_5_io_address),
    .io_dataRead(spriteMemories_5_io_dataRead)
  );
  Memory_73 spriteMemories_6 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_6_clock),
    .io_address(spriteMemories_6_io_address),
    .io_dataRead(spriteMemories_6_io_dataRead)
  );
  Memory_74 spriteMemories_7 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_7_clock),
    .io_address(spriteMemories_7_io_address),
    .io_dataRead(spriteMemories_7_io_dataRead)
  );
  Memory_75 spriteMemories_8 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_8_clock),
    .io_address(spriteMemories_8_io_address),
    .io_dataRead(spriteMemories_8_io_dataRead)
  );
  Memory_76 spriteMemories_9 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_9_clock),
    .io_address(spriteMemories_9_io_address),
    .io_dataRead(spriteMemories_9_io_dataRead)
  );
  Memory_77 spriteMemories_10 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_10_clock),
    .io_address(spriteMemories_10_io_address),
    .io_dataRead(spriteMemories_10_io_dataRead)
  );
  Memory_78 spriteMemories_11 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_11_clock),
    .io_address(spriteMemories_11_io_address),
    .io_dataRead(spriteMemories_11_io_dataRead)
  );
  Memory_79 spriteMemories_12 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_12_clock),
    .io_address(spriteMemories_12_io_address),
    .io_dataRead(spriteMemories_12_io_dataRead)
  );
  Memory_80 spriteMemories_13 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_13_clock),
    .io_address(spriteMemories_13_io_address),
    .io_dataRead(spriteMemories_13_io_dataRead)
  );
  Memory_81 spriteMemories_14 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_14_clock),
    .io_address(spriteMemories_14_io_address),
    .io_dataRead(spriteMemories_14_io_dataRead)
  );
  Memory_82 spriteMemories_15 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_15_clock),
    .io_address(spriteMemories_15_io_address),
    .io_dataRead(spriteMemories_15_io_dataRead)
  );
  Memory_83 spriteMemories_16 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_16_clock),
    .io_address(spriteMemories_16_io_address),
    .io_dataRead(spriteMemories_16_io_dataRead)
  );
  Memory_84 spriteMemories_17 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_17_clock),
    .io_address(spriteMemories_17_io_address),
    .io_dataRead(spriteMemories_17_io_dataRead)
  );
  Memory_85 spriteMemories_18 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_18_clock),
    .io_address(spriteMemories_18_io_address),
    .io_dataRead(spriteMemories_18_io_dataRead)
  );
  Memory_86 spriteMemories_19 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_19_clock),
    .io_address(spriteMemories_19_io_address),
    .io_dataRead(spriteMemories_19_io_dataRead)
  );
  Memory_87 spriteMemories_20 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_20_clock),
    .io_address(spriteMemories_20_io_address),
    .io_dataRead(spriteMemories_20_io_dataRead)
  );
  Memory_88 spriteMemories_21 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_21_clock),
    .io_address(spriteMemories_21_io_address),
    .io_dataRead(spriteMemories_21_io_dataRead)
  );
  Memory_89 spriteMemories_22 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_22_clock),
    .io_address(spriteMemories_22_io_address),
    .io_dataRead(spriteMemories_22_io_dataRead)
  );
  Memory_90 spriteMemories_23 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_23_clock),
    .io_address(spriteMemories_23_io_address),
    .io_dataRead(spriteMemories_23_io_dataRead)
  );
  Memory_91 spriteMemories_24 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_24_clock),
    .io_address(spriteMemories_24_io_address),
    .io_dataRead(spriteMemories_24_io_dataRead)
  );
  Memory_92 spriteMemories_25 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_25_clock),
    .io_address(spriteMemories_25_io_address),
    .io_dataRead(spriteMemories_25_io_dataRead)
  );
  Memory_93 spriteMemories_26 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_26_clock),
    .io_address(spriteMemories_26_io_address),
    .io_dataRead(spriteMemories_26_io_dataRead)
  );
  Memory_94 spriteMemories_27 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_27_clock),
    .io_address(spriteMemories_27_io_address),
    .io_dataRead(spriteMemories_27_io_dataRead)
  );
  Memory_95 spriteMemories_28 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_28_clock),
    .io_address(spriteMemories_28_io_address),
    .io_dataRead(spriteMemories_28_io_dataRead)
  );
  Memory_96 spriteMemories_29 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_29_clock),
    .io_address(spriteMemories_29_io_address),
    .io_dataRead(spriteMemories_29_io_dataRead)
  );
  Memory_97 spriteMemories_30 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_30_clock),
    .io_address(spriteMemories_30_io_address),
    .io_dataRead(spriteMemories_30_io_dataRead)
  );
  Memory_98 spriteMemories_31 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_31_clock),
    .io_address(spriteMemories_31_io_address),
    .io_dataRead(spriteMemories_31_io_dataRead)
  );
  Memory_99 spriteMemories_32 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_32_clock),
    .io_address(spriteMemories_32_io_address),
    .io_dataRead(spriteMemories_32_io_dataRead)
  );
  Memory_100 spriteMemories_33 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_33_clock),
    .io_address(spriteMemories_33_io_address),
    .io_dataRead(spriteMemories_33_io_dataRead)
  );
  Memory_101 spriteMemories_34 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_34_clock),
    .io_address(spriteMemories_34_io_address),
    .io_dataRead(spriteMemories_34_io_dataRead)
  );
  Memory_102 spriteMemories_35 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_35_clock),
    .io_address(spriteMemories_35_io_address),
    .io_dataRead(spriteMemories_35_io_dataRead)
  );
  Memory_103 spriteMemories_36 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_36_clock),
    .io_address(spriteMemories_36_io_address),
    .io_dataRead(spriteMemories_36_io_dataRead)
  );
  Memory_104 spriteMemories_37 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_37_clock),
    .io_address(spriteMemories_37_io_address),
    .io_dataRead(spriteMemories_37_io_dataRead)
  );
  Memory_105 spriteMemories_38 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_38_clock),
    .io_address(spriteMemories_38_io_address),
    .io_dataRead(spriteMemories_38_io_dataRead)
  );
  Memory_106 spriteMemories_39 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_39_clock),
    .io_address(spriteMemories_39_io_address),
    .io_dataRead(spriteMemories_39_io_dataRead)
  );
  Memory_107 spriteMemories_40 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_40_clock),
    .io_address(spriteMemories_40_io_address),
    .io_dataRead(spriteMemories_40_io_dataRead)
  );
  Memory_108 spriteMemories_41 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_41_clock),
    .io_address(spriteMemories_41_io_address),
    .io_dataRead(spriteMemories_41_io_dataRead)
  );
  Memory_109 spriteMemories_42 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_42_clock),
    .io_address(spriteMemories_42_io_address),
    .io_dataRead(spriteMemories_42_io_dataRead)
  );
  Memory_110 spriteMemories_43 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_43_clock),
    .io_address(spriteMemories_43_io_address),
    .io_dataRead(spriteMemories_43_io_dataRead)
  );
  Memory_111 spriteMemories_44 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_44_clock),
    .io_address(spriteMemories_44_io_address),
    .io_dataRead(spriteMemories_44_io_dataRead)
  );
  Memory_112 spriteMemories_45 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_45_clock),
    .io_address(spriteMemories_45_io_address),
    .io_dataRead(spriteMemories_45_io_dataRead)
  );
  Memory_113 spriteMemories_46 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_46_clock),
    .io_address(spriteMemories_46_io_address),
    .io_dataRead(spriteMemories_46_io_dataRead)
  );
  Memory_114 spriteMemories_47 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_47_clock),
    .io_address(spriteMemories_47_io_address),
    .io_dataRead(spriteMemories_47_io_dataRead)
  );
  Memory_115 spriteMemories_48 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_48_clock),
    .io_address(spriteMemories_48_io_address),
    .io_dataRead(spriteMemories_48_io_dataRead)
  );
  Memory_116 spriteMemories_49 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_49_clock),
    .io_address(spriteMemories_49_io_address),
    .io_dataRead(spriteMemories_49_io_dataRead)
  );
  Memory_117 spriteMemories_50 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_50_clock),
    .io_address(spriteMemories_50_io_address),
    .io_dataRead(spriteMemories_50_io_dataRead)
  );
  Memory_118 spriteMemories_51 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_51_clock),
    .io_address(spriteMemories_51_io_address),
    .io_dataRead(spriteMemories_51_io_dataRead)
  );
  Memory_119 spriteMemories_52 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_52_clock),
    .io_address(spriteMemories_52_io_address),
    .io_dataRead(spriteMemories_52_io_dataRead)
  );
  Memory_120 spriteMemories_53 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_53_clock),
    .io_address(spriteMemories_53_io_address),
    .io_dataRead(spriteMemories_53_io_dataRead)
  );
  Memory_121 spriteMemories_54 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_54_clock),
    .io_address(spriteMemories_54_io_address),
    .io_dataRead(spriteMemories_54_io_dataRead)
  );
  Memory_122 spriteMemories_55 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_55_clock),
    .io_address(spriteMemories_55_io_address),
    .io_dataRead(spriteMemories_55_io_dataRead)
  );
  Memory_123 spriteMemories_56 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_56_clock),
    .io_address(spriteMemories_56_io_address),
    .io_dataRead(spriteMemories_56_io_dataRead)
  );
  Memory_124 spriteMemories_57 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_57_clock),
    .io_address(spriteMemories_57_io_address),
    .io_dataRead(spriteMemories_57_io_dataRead)
  );
  Memory_125 spriteMemories_58 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_58_clock),
    .io_address(spriteMemories_58_io_address),
    .io_dataRead(spriteMemories_58_io_dataRead)
  );
  Memory_126 spriteMemories_59 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_59_clock),
    .io_address(spriteMemories_59_io_address),
    .io_dataRead(spriteMemories_59_io_dataRead)
  );
  Memory_127 spriteMemories_60 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_60_clock),
    .io_address(spriteMemories_60_io_address),
    .io_dataRead(spriteMemories_60_io_dataRead)
  );
  Memory_128 spriteMemories_61 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_61_clock),
    .io_address(spriteMemories_61_io_address),
    .io_dataRead(spriteMemories_61_io_dataRead)
  );
  Memory_129 spriteMemories_62 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_62_clock),
    .io_address(spriteMemories_62_io_address),
    .io_dataRead(spriteMemories_62_io_dataRead)
  );
  Memory_130 spriteMemories_63 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_63_clock),
    .io_address(spriteMemories_63_io_address),
    .io_dataRead(spriteMemories_63_io_dataRead)
  );
  Memory_131 spriteMemories_64 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_64_clock),
    .io_address(spriteMemories_64_io_address),
    .io_dataRead(spriteMemories_64_io_dataRead)
  );
  Memory_132 spriteMemories_65 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_65_clock),
    .io_address(spriteMemories_65_io_address),
    .io_dataRead(spriteMemories_65_io_dataRead)
  );
  Memory_133 spriteMemories_66 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_66_clock),
    .io_address(spriteMemories_66_io_address),
    .io_dataRead(spriteMemories_66_io_dataRead)
  );
  Memory_134 spriteMemories_67 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_67_clock),
    .io_address(spriteMemories_67_io_address),
    .io_dataRead(spriteMemories_67_io_dataRead)
  );
  Memory_135 spriteMemories_68 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_68_clock),
    .io_address(spriteMemories_68_io_address),
    .io_dataRead(spriteMemories_68_io_dataRead)
  );
  Memory_136 spriteMemories_69 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_69_clock),
    .io_address(spriteMemories_69_io_address),
    .io_dataRead(spriteMemories_69_io_dataRead)
  );
  Memory_137 spriteMemories_70 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_70_clock),
    .io_address(spriteMemories_70_io_address),
    .io_dataRead(spriteMemories_70_io_dataRead)
  );
  Memory_138 spriteMemories_71 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_71_clock),
    .io_address(spriteMemories_71_io_address),
    .io_dataRead(spriteMemories_71_io_dataRead)
  );
  Memory_139 spriteMemories_72 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_72_clock),
    .io_address(spriteMemories_72_io_address),
    .io_dataRead(spriteMemories_72_io_dataRead)
  );
  Memory_140 spriteMemories_73 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_73_clock),
    .io_address(spriteMemories_73_io_address),
    .io_dataRead(spriteMemories_73_io_dataRead)
  );
  Memory_141 spriteMemories_74 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_74_clock),
    .io_address(spriteMemories_74_io_address),
    .io_dataRead(spriteMemories_74_io_dataRead)
  );
  Memory_142 spriteMemories_75 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_75_clock),
    .io_address(spriteMemories_75_io_address),
    .io_dataRead(spriteMemories_75_io_dataRead)
  );
  Memory_143 spriteMemories_76 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_76_clock),
    .io_address(spriteMemories_76_io_address),
    .io_dataRead(spriteMemories_76_io_dataRead)
  );
  Memory_144 spriteMemories_77 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_77_clock),
    .io_address(spriteMemories_77_io_address),
    .io_dataRead(spriteMemories_77_io_dataRead)
  );
  Memory_145 spriteMemories_78 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_78_clock),
    .io_address(spriteMemories_78_io_address),
    .io_dataRead(spriteMemories_78_io_dataRead)
  );
  Memory_146 spriteMemories_79 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_79_clock),
    .io_address(spriteMemories_79_io_address),
    .io_dataRead(spriteMemories_79_io_dataRead)
  );
  Memory_147 spriteMemories_80 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_80_clock),
    .io_address(spriteMemories_80_io_address),
    .io_dataRead(spriteMemories_80_io_dataRead)
  );
  Memory_148 spriteMemories_81 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_81_clock),
    .io_address(spriteMemories_81_io_address),
    .io_dataRead(spriteMemories_81_io_dataRead)
  );
  Memory_149 spriteMemories_82 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_82_clock),
    .io_address(spriteMemories_82_io_address),
    .io_dataRead(spriteMemories_82_io_dataRead)
  );
  Memory_150 spriteMemories_83 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_83_clock),
    .io_address(spriteMemories_83_io_address),
    .io_dataRead(spriteMemories_83_io_dataRead)
  );
  Memory_151 spriteMemories_84 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_84_clock),
    .io_address(spriteMemories_84_io_address),
    .io_dataRead(spriteMemories_84_io_dataRead)
  );
  Memory_152 spriteMemories_85 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_85_clock),
    .io_address(spriteMemories_85_io_address),
    .io_dataRead(spriteMemories_85_io_dataRead)
  );
  Memory_153 spriteMemories_86 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_86_clock),
    .io_address(spriteMemories_86_io_address),
    .io_dataRead(spriteMemories_86_io_dataRead)
  );
  Memory_154 spriteMemories_87 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_87_clock),
    .io_address(spriteMemories_87_io_address),
    .io_dataRead(spriteMemories_87_io_dataRead)
  );
  Memory_155 spriteMemories_88 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_88_clock),
    .io_address(spriteMemories_88_io_address),
    .io_dataRead(spriteMemories_88_io_dataRead)
  );
  Memory_156 spriteMemories_89 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_89_clock),
    .io_address(spriteMemories_89_io_address),
    .io_dataRead(spriteMemories_89_io_dataRead)
  );
  Memory_157 spriteMemories_90 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_90_clock),
    .io_address(spriteMemories_90_io_address),
    .io_dataRead(spriteMemories_90_io_dataRead)
  );
  Memory_158 spriteMemories_91 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_91_clock),
    .io_address(spriteMemories_91_io_address),
    .io_dataRead(spriteMemories_91_io_dataRead)
  );
  Memory_159 spriteMemories_92 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_92_clock),
    .io_address(spriteMemories_92_io_address),
    .io_dataRead(spriteMemories_92_io_dataRead)
  );
  Memory_160 spriteMemories_93 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_93_clock),
    .io_address(spriteMemories_93_io_address),
    .io_dataRead(spriteMemories_93_io_dataRead)
  );
  Memory_161 spriteMemories_94 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_94_clock),
    .io_address(spriteMemories_94_io_address),
    .io_dataRead(spriteMemories_94_io_dataRead)
  );
  Memory_162 spriteMemories_95 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_95_clock),
    .io_address(spriteMemories_95_io_address),
    .io_dataRead(spriteMemories_95_io_dataRead)
  );
  Memory_163 spriteMemories_96 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_96_clock),
    .io_address(spriteMemories_96_io_address),
    .io_dataRead(spriteMemories_96_io_dataRead)
  );
  Memory_164 spriteMemories_97 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_97_clock),
    .io_address(spriteMemories_97_io_address),
    .io_dataRead(spriteMemories_97_io_dataRead)
  );
  Memory_165 spriteMemories_98 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_98_clock),
    .io_address(spriteMemories_98_io_address),
    .io_dataRead(spriteMemories_98_io_dataRead)
  );
  Memory_166 spriteMemories_99 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_99_clock),
    .io_address(spriteMemories_99_io_address),
    .io_dataRead(spriteMemories_99_io_dataRead)
  );
  Memory_167 spriteMemories_100 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_100_clock),
    .io_address(spriteMemories_100_io_address),
    .io_dataRead(spriteMemories_100_io_dataRead)
  );
  Memory_168 spriteMemories_101 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_101_clock),
    .io_address(spriteMemories_101_io_address),
    .io_dataRead(spriteMemories_101_io_dataRead)
  );
  Memory_169 spriteMemories_102 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_102_clock),
    .io_address(spriteMemories_102_io_address),
    .io_dataRead(spriteMemories_102_io_dataRead)
  );
  Memory_170 spriteMemories_103 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_103_clock),
    .io_address(spriteMemories_103_io_address),
    .io_dataRead(spriteMemories_103_io_dataRead)
  );
  Memory_171 spriteMemories_104 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_104_clock),
    .io_address(spriteMemories_104_io_address),
    .io_dataRead(spriteMemories_104_io_dataRead)
  );
  Memory_172 spriteMemories_105 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_105_clock),
    .io_address(spriteMemories_105_io_address),
    .io_dataRead(spriteMemories_105_io_dataRead)
  );
  Memory_173 spriteMemories_106 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_106_clock),
    .io_address(spriteMemories_106_io_address),
    .io_dataRead(spriteMemories_106_io_dataRead)
  );
  Memory_174 spriteMemories_107 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_107_clock),
    .io_address(spriteMemories_107_io_address),
    .io_dataRead(spriteMemories_107_io_dataRead)
  );
  Memory_175 spriteMemories_108 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_108_clock),
    .io_address(spriteMemories_108_io_address),
    .io_dataRead(spriteMemories_108_io_dataRead)
  );
  Memory_176 spriteMemories_109 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_109_clock),
    .io_address(spriteMemories_109_io_address),
    .io_dataRead(spriteMemories_109_io_dataRead)
  );
  Memory_177 spriteMemories_110 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_110_clock),
    .io_address(spriteMemories_110_io_address),
    .io_dataRead(spriteMemories_110_io_dataRead)
  );
  Memory_178 spriteMemories_111 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_111_clock),
    .io_address(spriteMemories_111_io_address),
    .io_dataRead(spriteMemories_111_io_dataRead)
  );
  Memory_179 spriteMemories_112 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_112_clock),
    .io_address(spriteMemories_112_io_address),
    .io_dataRead(spriteMemories_112_io_dataRead)
  );
  Memory_180 spriteMemories_113 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_113_clock),
    .io_address(spriteMemories_113_io_address),
    .io_dataRead(spriteMemories_113_io_dataRead)
  );
  Memory_181 spriteMemories_114 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_114_clock),
    .io_address(spriteMemories_114_io_address),
    .io_dataRead(spriteMemories_114_io_dataRead)
  );
  Memory_182 spriteMemories_115 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_115_clock),
    .io_address(spriteMemories_115_io_address),
    .io_dataRead(spriteMemories_115_io_dataRead)
  );
  Memory_183 spriteMemories_116 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_116_clock),
    .io_address(spriteMemories_116_io_address),
    .io_dataRead(spriteMemories_116_io_dataRead)
  );
  Memory_184 spriteMemories_117 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_117_clock),
    .io_address(spriteMemories_117_io_address),
    .io_dataRead(spriteMemories_117_io_dataRead)
  );
  Memory_185 spriteMemories_118 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_118_clock),
    .io_address(spriteMemories_118_io_address),
    .io_dataRead(spriteMemories_118_io_dataRead)
  );
  Memory_186 spriteMemories_119 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_119_clock),
    .io_address(spriteMemories_119_io_address),
    .io_dataRead(spriteMemories_119_io_dataRead)
  );
  Memory_187 spriteMemories_120 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_120_clock),
    .io_address(spriteMemories_120_io_address),
    .io_dataRead(spriteMemories_120_io_dataRead)
  );
  Memory_188 spriteMemories_121 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_121_clock),
    .io_address(spriteMemories_121_io_address),
    .io_dataRead(spriteMemories_121_io_dataRead)
  );
  Memory_189 spriteMemories_122 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_122_clock),
    .io_address(spriteMemories_122_io_address),
    .io_dataRead(spriteMemories_122_io_dataRead)
  );
  Memory_190 spriteMemories_123 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_123_clock),
    .io_address(spriteMemories_123_io_address),
    .io_dataRead(spriteMemories_123_io_dataRead)
  );
  Memory_191 spriteMemories_124 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_124_clock),
    .io_address(spriteMemories_124_io_address),
    .io_dataRead(spriteMemories_124_io_dataRead)
  );
  Memory_192 spriteMemories_125 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_125_clock),
    .io_address(spriteMemories_125_io_address),
    .io_dataRead(spriteMemories_125_io_dataRead)
  );
  Memory_193 spriteMemories_126 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_126_clock),
    .io_address(spriteMemories_126_io_address),
    .io_dataRead(spriteMemories_126_io_dataRead)
  );
  Memory_194 spriteMemories_127 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_127_clock),
    .io_address(spriteMemories_127_io_address),
    .io_dataRead(spriteMemories_127_io_dataRead)
  );
  MultiHotPriortyReductionTree multiHotPriortyReductionTree ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
    .io_dataInput_0(multiHotPriortyReductionTree_io_dataInput_0),
    .io_dataInput_1(multiHotPriortyReductionTree_io_dataInput_1),
    .io_dataInput_2(multiHotPriortyReductionTree_io_dataInput_2),
    .io_dataInput_3(multiHotPriortyReductionTree_io_dataInput_3),
    .io_dataInput_4(multiHotPriortyReductionTree_io_dataInput_4),
    .io_dataInput_5(multiHotPriortyReductionTree_io_dataInput_5),
    .io_dataInput_6(multiHotPriortyReductionTree_io_dataInput_6),
    .io_dataInput_7(multiHotPriortyReductionTree_io_dataInput_7),
    .io_dataInput_8(multiHotPriortyReductionTree_io_dataInput_8),
    .io_dataInput_9(multiHotPriortyReductionTree_io_dataInput_9),
    .io_dataInput_10(multiHotPriortyReductionTree_io_dataInput_10),
    .io_dataInput_11(multiHotPriortyReductionTree_io_dataInput_11),
    .io_dataInput_12(multiHotPriortyReductionTree_io_dataInput_12),
    .io_dataInput_13(multiHotPriortyReductionTree_io_dataInput_13),
    .io_dataInput_14(multiHotPriortyReductionTree_io_dataInput_14),
    .io_dataInput_15(multiHotPriortyReductionTree_io_dataInput_15),
    .io_dataInput_16(multiHotPriortyReductionTree_io_dataInput_16),
    .io_dataInput_17(multiHotPriortyReductionTree_io_dataInput_17),
    .io_dataInput_18(multiHotPriortyReductionTree_io_dataInput_18),
    .io_dataInput_19(multiHotPriortyReductionTree_io_dataInput_19),
    .io_dataInput_20(multiHotPriortyReductionTree_io_dataInput_20),
    .io_dataInput_21(multiHotPriortyReductionTree_io_dataInput_21),
    .io_dataInput_22(multiHotPriortyReductionTree_io_dataInput_22),
    .io_dataInput_23(multiHotPriortyReductionTree_io_dataInput_23),
    .io_dataInput_24(multiHotPriortyReductionTree_io_dataInput_24),
    .io_dataInput_25(multiHotPriortyReductionTree_io_dataInput_25),
    .io_dataInput_26(multiHotPriortyReductionTree_io_dataInput_26),
    .io_dataInput_27(multiHotPriortyReductionTree_io_dataInput_27),
    .io_dataInput_28(multiHotPriortyReductionTree_io_dataInput_28),
    .io_dataInput_29(multiHotPriortyReductionTree_io_dataInput_29),
    .io_dataInput_30(multiHotPriortyReductionTree_io_dataInput_30),
    .io_dataInput_31(multiHotPriortyReductionTree_io_dataInput_31),
    .io_dataInput_32(multiHotPriortyReductionTree_io_dataInput_32),
    .io_dataInput_33(multiHotPriortyReductionTree_io_dataInput_33),
    .io_dataInput_34(multiHotPriortyReductionTree_io_dataInput_34),
    .io_dataInput_35(multiHotPriortyReductionTree_io_dataInput_35),
    .io_dataInput_36(multiHotPriortyReductionTree_io_dataInput_36),
    .io_dataInput_37(multiHotPriortyReductionTree_io_dataInput_37),
    .io_dataInput_38(multiHotPriortyReductionTree_io_dataInput_38),
    .io_dataInput_39(multiHotPriortyReductionTree_io_dataInput_39),
    .io_dataInput_40(multiHotPriortyReductionTree_io_dataInput_40),
    .io_dataInput_41(multiHotPriortyReductionTree_io_dataInput_41),
    .io_dataInput_42(multiHotPriortyReductionTree_io_dataInput_42),
    .io_dataInput_43(multiHotPriortyReductionTree_io_dataInput_43),
    .io_dataInput_44(multiHotPriortyReductionTree_io_dataInput_44),
    .io_dataInput_45(multiHotPriortyReductionTree_io_dataInput_45),
    .io_dataInput_46(multiHotPriortyReductionTree_io_dataInput_46),
    .io_dataInput_47(multiHotPriortyReductionTree_io_dataInput_47),
    .io_dataInput_48(multiHotPriortyReductionTree_io_dataInput_48),
    .io_dataInput_49(multiHotPriortyReductionTree_io_dataInput_49),
    .io_dataInput_50(multiHotPriortyReductionTree_io_dataInput_50),
    .io_dataInput_51(multiHotPriortyReductionTree_io_dataInput_51),
    .io_dataInput_52(multiHotPriortyReductionTree_io_dataInput_52),
    .io_dataInput_53(multiHotPriortyReductionTree_io_dataInput_53),
    .io_dataInput_54(multiHotPriortyReductionTree_io_dataInput_54),
    .io_dataInput_55(multiHotPriortyReductionTree_io_dataInput_55),
    .io_dataInput_56(multiHotPriortyReductionTree_io_dataInput_56),
    .io_dataInput_57(multiHotPriortyReductionTree_io_dataInput_57),
    .io_dataInput_58(multiHotPriortyReductionTree_io_dataInput_58),
    .io_dataInput_59(multiHotPriortyReductionTree_io_dataInput_59),
    .io_dataInput_60(multiHotPriortyReductionTree_io_dataInput_60),
    .io_dataInput_61(multiHotPriortyReductionTree_io_dataInput_61),
    .io_dataInput_62(multiHotPriortyReductionTree_io_dataInput_62),
    .io_dataInput_63(multiHotPriortyReductionTree_io_dataInput_63),
    .io_dataInput_64(multiHotPriortyReductionTree_io_dataInput_64),
    .io_dataInput_65(multiHotPriortyReductionTree_io_dataInput_65),
    .io_dataInput_66(multiHotPriortyReductionTree_io_dataInput_66),
    .io_dataInput_67(multiHotPriortyReductionTree_io_dataInput_67),
    .io_dataInput_68(multiHotPriortyReductionTree_io_dataInput_68),
    .io_dataInput_69(multiHotPriortyReductionTree_io_dataInput_69),
    .io_dataInput_70(multiHotPriortyReductionTree_io_dataInput_70),
    .io_dataInput_71(multiHotPriortyReductionTree_io_dataInput_71),
    .io_dataInput_72(multiHotPriortyReductionTree_io_dataInput_72),
    .io_dataInput_73(multiHotPriortyReductionTree_io_dataInput_73),
    .io_dataInput_74(multiHotPriortyReductionTree_io_dataInput_74),
    .io_dataInput_75(multiHotPriortyReductionTree_io_dataInput_75),
    .io_dataInput_76(multiHotPriortyReductionTree_io_dataInput_76),
    .io_dataInput_77(multiHotPriortyReductionTree_io_dataInput_77),
    .io_dataInput_78(multiHotPriortyReductionTree_io_dataInput_78),
    .io_dataInput_79(multiHotPriortyReductionTree_io_dataInput_79),
    .io_dataInput_80(multiHotPriortyReductionTree_io_dataInput_80),
    .io_dataInput_81(multiHotPriortyReductionTree_io_dataInput_81),
    .io_dataInput_82(multiHotPriortyReductionTree_io_dataInput_82),
    .io_dataInput_83(multiHotPriortyReductionTree_io_dataInput_83),
    .io_dataInput_84(multiHotPriortyReductionTree_io_dataInput_84),
    .io_dataInput_85(multiHotPriortyReductionTree_io_dataInput_85),
    .io_dataInput_86(multiHotPriortyReductionTree_io_dataInput_86),
    .io_dataInput_87(multiHotPriortyReductionTree_io_dataInput_87),
    .io_dataInput_88(multiHotPriortyReductionTree_io_dataInput_88),
    .io_dataInput_89(multiHotPriortyReductionTree_io_dataInput_89),
    .io_dataInput_90(multiHotPriortyReductionTree_io_dataInput_90),
    .io_dataInput_91(multiHotPriortyReductionTree_io_dataInput_91),
    .io_dataInput_92(multiHotPriortyReductionTree_io_dataInput_92),
    .io_dataInput_93(multiHotPriortyReductionTree_io_dataInput_93),
    .io_dataInput_94(multiHotPriortyReductionTree_io_dataInput_94),
    .io_dataInput_95(multiHotPriortyReductionTree_io_dataInput_95),
    .io_dataInput_96(multiHotPriortyReductionTree_io_dataInput_96),
    .io_dataInput_97(multiHotPriortyReductionTree_io_dataInput_97),
    .io_dataInput_98(multiHotPriortyReductionTree_io_dataInput_98),
    .io_dataInput_99(multiHotPriortyReductionTree_io_dataInput_99),
    .io_dataInput_100(multiHotPriortyReductionTree_io_dataInput_100),
    .io_dataInput_101(multiHotPriortyReductionTree_io_dataInput_101),
    .io_dataInput_102(multiHotPriortyReductionTree_io_dataInput_102),
    .io_dataInput_103(multiHotPriortyReductionTree_io_dataInput_103),
    .io_dataInput_104(multiHotPriortyReductionTree_io_dataInput_104),
    .io_dataInput_105(multiHotPriortyReductionTree_io_dataInput_105),
    .io_dataInput_106(multiHotPriortyReductionTree_io_dataInput_106),
    .io_dataInput_107(multiHotPriortyReductionTree_io_dataInput_107),
    .io_dataInput_108(multiHotPriortyReductionTree_io_dataInput_108),
    .io_dataInput_109(multiHotPriortyReductionTree_io_dataInput_109),
    .io_dataInput_110(multiHotPriortyReductionTree_io_dataInput_110),
    .io_dataInput_111(multiHotPriortyReductionTree_io_dataInput_111),
    .io_dataInput_112(multiHotPriortyReductionTree_io_dataInput_112),
    .io_dataInput_113(multiHotPriortyReductionTree_io_dataInput_113),
    .io_dataInput_114(multiHotPriortyReductionTree_io_dataInput_114),
    .io_dataInput_115(multiHotPriortyReductionTree_io_dataInput_115),
    .io_dataInput_116(multiHotPriortyReductionTree_io_dataInput_116),
    .io_dataInput_117(multiHotPriortyReductionTree_io_dataInput_117),
    .io_dataInput_118(multiHotPriortyReductionTree_io_dataInput_118),
    .io_dataInput_119(multiHotPriortyReductionTree_io_dataInput_119),
    .io_dataInput_120(multiHotPriortyReductionTree_io_dataInput_120),
    .io_dataInput_121(multiHotPriortyReductionTree_io_dataInput_121),
    .io_dataInput_122(multiHotPriortyReductionTree_io_dataInput_122),
    .io_dataInput_123(multiHotPriortyReductionTree_io_dataInput_123),
    .io_dataInput_124(multiHotPriortyReductionTree_io_dataInput_124),
    .io_dataInput_125(multiHotPriortyReductionTree_io_dataInput_125),
    .io_dataInput_126(multiHotPriortyReductionTree_io_dataInput_126),
    .io_dataInput_127(multiHotPriortyReductionTree_io_dataInput_127),
    .io_selectInput_0(multiHotPriortyReductionTree_io_selectInput_0),
    .io_selectInput_1(multiHotPriortyReductionTree_io_selectInput_1),
    .io_selectInput_2(multiHotPriortyReductionTree_io_selectInput_2),
    .io_selectInput_3(multiHotPriortyReductionTree_io_selectInput_3),
    .io_selectInput_4(multiHotPriortyReductionTree_io_selectInput_4),
    .io_selectInput_5(multiHotPriortyReductionTree_io_selectInput_5),
    .io_selectInput_6(multiHotPriortyReductionTree_io_selectInput_6),
    .io_selectInput_7(multiHotPriortyReductionTree_io_selectInput_7),
    .io_selectInput_8(multiHotPriortyReductionTree_io_selectInput_8),
    .io_selectInput_9(multiHotPriortyReductionTree_io_selectInput_9),
    .io_selectInput_10(multiHotPriortyReductionTree_io_selectInput_10),
    .io_selectInput_11(multiHotPriortyReductionTree_io_selectInput_11),
    .io_selectInput_12(multiHotPriortyReductionTree_io_selectInput_12),
    .io_selectInput_13(multiHotPriortyReductionTree_io_selectInput_13),
    .io_selectInput_14(multiHotPriortyReductionTree_io_selectInput_14),
    .io_selectInput_15(multiHotPriortyReductionTree_io_selectInput_15),
    .io_selectInput_16(multiHotPriortyReductionTree_io_selectInput_16),
    .io_selectInput_17(multiHotPriortyReductionTree_io_selectInput_17),
    .io_selectInput_18(multiHotPriortyReductionTree_io_selectInput_18),
    .io_selectInput_19(multiHotPriortyReductionTree_io_selectInput_19),
    .io_selectInput_20(multiHotPriortyReductionTree_io_selectInput_20),
    .io_selectInput_21(multiHotPriortyReductionTree_io_selectInput_21),
    .io_selectInput_22(multiHotPriortyReductionTree_io_selectInput_22),
    .io_selectInput_23(multiHotPriortyReductionTree_io_selectInput_23),
    .io_selectInput_24(multiHotPriortyReductionTree_io_selectInput_24),
    .io_selectInput_25(multiHotPriortyReductionTree_io_selectInput_25),
    .io_selectInput_26(multiHotPriortyReductionTree_io_selectInput_26),
    .io_selectInput_27(multiHotPriortyReductionTree_io_selectInput_27),
    .io_selectInput_28(multiHotPriortyReductionTree_io_selectInput_28),
    .io_selectInput_29(multiHotPriortyReductionTree_io_selectInput_29),
    .io_selectInput_30(multiHotPriortyReductionTree_io_selectInput_30),
    .io_selectInput_31(multiHotPriortyReductionTree_io_selectInput_31),
    .io_selectInput_32(multiHotPriortyReductionTree_io_selectInput_32),
    .io_selectInput_33(multiHotPriortyReductionTree_io_selectInput_33),
    .io_selectInput_34(multiHotPriortyReductionTree_io_selectInput_34),
    .io_selectInput_35(multiHotPriortyReductionTree_io_selectInput_35),
    .io_selectInput_36(multiHotPriortyReductionTree_io_selectInput_36),
    .io_selectInput_37(multiHotPriortyReductionTree_io_selectInput_37),
    .io_selectInput_38(multiHotPriortyReductionTree_io_selectInput_38),
    .io_selectInput_39(multiHotPriortyReductionTree_io_selectInput_39),
    .io_selectInput_40(multiHotPriortyReductionTree_io_selectInput_40),
    .io_selectInput_41(multiHotPriortyReductionTree_io_selectInput_41),
    .io_selectInput_42(multiHotPriortyReductionTree_io_selectInput_42),
    .io_selectInput_43(multiHotPriortyReductionTree_io_selectInput_43),
    .io_selectInput_44(multiHotPriortyReductionTree_io_selectInput_44),
    .io_selectInput_45(multiHotPriortyReductionTree_io_selectInput_45),
    .io_selectInput_46(multiHotPriortyReductionTree_io_selectInput_46),
    .io_selectInput_47(multiHotPriortyReductionTree_io_selectInput_47),
    .io_selectInput_48(multiHotPriortyReductionTree_io_selectInput_48),
    .io_selectInput_49(multiHotPriortyReductionTree_io_selectInput_49),
    .io_selectInput_50(multiHotPriortyReductionTree_io_selectInput_50),
    .io_selectInput_51(multiHotPriortyReductionTree_io_selectInput_51),
    .io_selectInput_52(multiHotPriortyReductionTree_io_selectInput_52),
    .io_selectInput_53(multiHotPriortyReductionTree_io_selectInput_53),
    .io_selectInput_54(multiHotPriortyReductionTree_io_selectInput_54),
    .io_selectInput_55(multiHotPriortyReductionTree_io_selectInput_55),
    .io_selectInput_56(multiHotPriortyReductionTree_io_selectInput_56),
    .io_selectInput_57(multiHotPriortyReductionTree_io_selectInput_57),
    .io_selectInput_58(multiHotPriortyReductionTree_io_selectInput_58),
    .io_selectInput_59(multiHotPriortyReductionTree_io_selectInput_59),
    .io_selectInput_60(multiHotPriortyReductionTree_io_selectInput_60),
    .io_selectInput_61(multiHotPriortyReductionTree_io_selectInput_61),
    .io_selectInput_62(multiHotPriortyReductionTree_io_selectInput_62),
    .io_selectInput_63(multiHotPriortyReductionTree_io_selectInput_63),
    .io_selectInput_64(multiHotPriortyReductionTree_io_selectInput_64),
    .io_selectInput_65(multiHotPriortyReductionTree_io_selectInput_65),
    .io_selectInput_66(multiHotPriortyReductionTree_io_selectInput_66),
    .io_selectInput_67(multiHotPriortyReductionTree_io_selectInput_67),
    .io_selectInput_68(multiHotPriortyReductionTree_io_selectInput_68),
    .io_selectInput_69(multiHotPriortyReductionTree_io_selectInput_69),
    .io_selectInput_70(multiHotPriortyReductionTree_io_selectInput_70),
    .io_selectInput_71(multiHotPriortyReductionTree_io_selectInput_71),
    .io_selectInput_72(multiHotPriortyReductionTree_io_selectInput_72),
    .io_selectInput_73(multiHotPriortyReductionTree_io_selectInput_73),
    .io_selectInput_74(multiHotPriortyReductionTree_io_selectInput_74),
    .io_selectInput_75(multiHotPriortyReductionTree_io_selectInput_75),
    .io_selectInput_76(multiHotPriortyReductionTree_io_selectInput_76),
    .io_selectInput_77(multiHotPriortyReductionTree_io_selectInput_77),
    .io_selectInput_78(multiHotPriortyReductionTree_io_selectInput_78),
    .io_selectInput_79(multiHotPriortyReductionTree_io_selectInput_79),
    .io_selectInput_80(multiHotPriortyReductionTree_io_selectInput_80),
    .io_selectInput_81(multiHotPriortyReductionTree_io_selectInput_81),
    .io_selectInput_82(multiHotPriortyReductionTree_io_selectInput_82),
    .io_selectInput_83(multiHotPriortyReductionTree_io_selectInput_83),
    .io_selectInput_84(multiHotPriortyReductionTree_io_selectInput_84),
    .io_selectInput_85(multiHotPriortyReductionTree_io_selectInput_85),
    .io_selectInput_86(multiHotPriortyReductionTree_io_selectInput_86),
    .io_selectInput_87(multiHotPriortyReductionTree_io_selectInput_87),
    .io_selectInput_88(multiHotPriortyReductionTree_io_selectInput_88),
    .io_selectInput_89(multiHotPriortyReductionTree_io_selectInput_89),
    .io_selectInput_90(multiHotPriortyReductionTree_io_selectInput_90),
    .io_selectInput_91(multiHotPriortyReductionTree_io_selectInput_91),
    .io_selectInput_92(multiHotPriortyReductionTree_io_selectInput_92),
    .io_selectInput_93(multiHotPriortyReductionTree_io_selectInput_93),
    .io_selectInput_94(multiHotPriortyReductionTree_io_selectInput_94),
    .io_selectInput_95(multiHotPriortyReductionTree_io_selectInput_95),
    .io_selectInput_96(multiHotPriortyReductionTree_io_selectInput_96),
    .io_selectInput_97(multiHotPriortyReductionTree_io_selectInput_97),
    .io_selectInput_98(multiHotPriortyReductionTree_io_selectInput_98),
    .io_selectInput_99(multiHotPriortyReductionTree_io_selectInput_99),
    .io_selectInput_100(multiHotPriortyReductionTree_io_selectInput_100),
    .io_selectInput_101(multiHotPriortyReductionTree_io_selectInput_101),
    .io_selectInput_102(multiHotPriortyReductionTree_io_selectInput_102),
    .io_selectInput_103(multiHotPriortyReductionTree_io_selectInput_103),
    .io_selectInput_104(multiHotPriortyReductionTree_io_selectInput_104),
    .io_selectInput_105(multiHotPriortyReductionTree_io_selectInput_105),
    .io_selectInput_106(multiHotPriortyReductionTree_io_selectInput_106),
    .io_selectInput_107(multiHotPriortyReductionTree_io_selectInput_107),
    .io_selectInput_108(multiHotPriortyReductionTree_io_selectInput_108),
    .io_selectInput_109(multiHotPriortyReductionTree_io_selectInput_109),
    .io_selectInput_110(multiHotPriortyReductionTree_io_selectInput_110),
    .io_selectInput_111(multiHotPriortyReductionTree_io_selectInput_111),
    .io_selectInput_112(multiHotPriortyReductionTree_io_selectInput_112),
    .io_selectInput_113(multiHotPriortyReductionTree_io_selectInput_113),
    .io_selectInput_114(multiHotPriortyReductionTree_io_selectInput_114),
    .io_selectInput_115(multiHotPriortyReductionTree_io_selectInput_115),
    .io_selectInput_116(multiHotPriortyReductionTree_io_selectInput_116),
    .io_selectInput_117(multiHotPriortyReductionTree_io_selectInput_117),
    .io_selectInput_118(multiHotPriortyReductionTree_io_selectInput_118),
    .io_selectInput_119(multiHotPriortyReductionTree_io_selectInput_119),
    .io_selectInput_120(multiHotPriortyReductionTree_io_selectInput_120),
    .io_selectInput_121(multiHotPriortyReductionTree_io_selectInput_121),
    .io_selectInput_122(multiHotPriortyReductionTree_io_selectInput_122),
    .io_selectInput_123(multiHotPriortyReductionTree_io_selectInput_123),
    .io_selectInput_124(multiHotPriortyReductionTree_io_selectInput_124),
    .io_selectInput_125(multiHotPriortyReductionTree_io_selectInput_125),
    .io_selectInput_126(multiHotPriortyReductionTree_io_selectInput_126),
    .io_selectInput_127(multiHotPriortyReductionTree_io_selectInput_127),
    .io_dataOutput(multiHotPriortyReductionTree_io_dataOutput),
    .io_selectOutput(multiHotPriortyReductionTree_io_selectOutput)
  );
  assign io_newFrame = run & _GEN_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13 71:15]
  assign io_missingFrameError = missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 131:24]
  assign io_viewBoxOutOfRangeError = viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 133:29]
  assign io_vgaRed = io_vgaRed_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 349:13]
  assign io_vgaBlue = io_vgaBlue_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 351:14]
  assign io_vgaGreen = io_vgaGreen_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 350:15]
  assign io_Hsync = io_Hsync_pipeReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 94:12]
  assign io_Vsync = io_Vsync_pipeReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 95:12]
  assign backTileMemories_0_clock = clock;
  assign backTileMemories_0_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_1_clock = clock;
  assign backTileMemories_1_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_2_clock = clock;
  assign backTileMemories_2_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_3_clock = clock;
  assign backTileMemories_3_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_4_clock = clock;
  assign backTileMemories_4_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_5_clock = clock;
  assign backTileMemories_5_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_6_clock = clock;
  assign backTileMemories_6_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_7_clock = clock;
  assign backTileMemories_7_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_8_clock = clock;
  assign backTileMemories_8_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_9_clock = clock;
  assign backTileMemories_9_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_10_clock = clock;
  assign backTileMemories_10_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_11_clock = clock;
  assign backTileMemories_11_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_12_clock = clock;
  assign backTileMemories_12_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_13_clock = clock;
  assign backTileMemories_13_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_14_clock = clock;
  assign backTileMemories_14_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_15_clock = clock;
  assign backTileMemories_15_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_16_clock = clock;
  assign backTileMemories_16_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_17_clock = clock;
  assign backTileMemories_17_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_18_clock = clock;
  assign backTileMemories_18_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_19_clock = clock;
  assign backTileMemories_19_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_20_clock = clock;
  assign backTileMemories_20_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_21_clock = clock;
  assign backTileMemories_21_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_22_clock = clock;
  assign backTileMemories_22_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_23_clock = clock;
  assign backTileMemories_23_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_24_clock = clock;
  assign backTileMemories_24_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_25_clock = clock;
  assign backTileMemories_25_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_26_clock = clock;
  assign backTileMemories_26_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_27_clock = clock;
  assign backTileMemories_27_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_28_clock = clock;
  assign backTileMemories_28_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_29_clock = clock;
  assign backTileMemories_29_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_30_clock = clock;
  assign backTileMemories_30_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_31_clock = clock;
  assign backTileMemories_31_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_32_clock = clock;
  assign backTileMemories_32_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_33_clock = clock;
  assign backTileMemories_33_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_34_clock = clock;
  assign backTileMemories_34_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_35_clock = clock;
  assign backTileMemories_35_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_36_clock = clock;
  assign backTileMemories_36_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_37_clock = clock;
  assign backTileMemories_37_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_38_clock = clock;
  assign backTileMemories_38_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_39_clock = clock;
  assign backTileMemories_39_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_40_clock = clock;
  assign backTileMemories_40_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_41_clock = clock;
  assign backTileMemories_41_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_42_clock = clock;
  assign backTileMemories_42_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_43_clock = clock;
  assign backTileMemories_43_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_44_clock = clock;
  assign backTileMemories_44_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_45_clock = clock;
  assign backTileMemories_45_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_46_clock = clock;
  assign backTileMemories_46_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_47_clock = clock;
  assign backTileMemories_47_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_48_clock = clock;
  assign backTileMemories_48_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_49_clock = clock;
  assign backTileMemories_49_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_50_clock = clock;
  assign backTileMemories_50_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_51_clock = clock;
  assign backTileMemories_51_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_52_clock = clock;
  assign backTileMemories_52_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_53_clock = clock;
  assign backTileMemories_53_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_54_clock = clock;
  assign backTileMemories_54_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_55_clock = clock;
  assign backTileMemories_55_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_56_clock = clock;
  assign backTileMemories_56_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_57_clock = clock;
  assign backTileMemories_57_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_58_clock = clock;
  assign backTileMemories_58_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_59_clock = clock;
  assign backTileMemories_59_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_60_clock = clock;
  assign backTileMemories_60_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_61_clock = clock;
  assign backTileMemories_61_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_62_clock = clock;
  assign backTileMemories_62_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_63_clock = clock;
  assign backTileMemories_63_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backBufferMemory_clock = clock;
  assign backBufferMemory_io_address = _backBufferMemory_io_address_T_5[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:31]
  assign backBufferMemory_io_writeEnable = copyEnabledReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 228:35]
  assign backBufferMemory_io_dataWrite = backBufferShadowMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 229:33]
  assign backBufferShadowMemory_clock = clock;
  assign backBufferShadowMemory_io_address = restoreEnabled ? backBufferShadowMemory_io_address_REG :
    _backBufferShadowMemory_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:43]
  assign backBufferShadowMemory_io_writeEnable = restoreEnabled & backBufferShadowMemory_io_writeEnable_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:47]
  assign backBufferShadowMemory_io_dataWrite = restoreEnabled ? backBufferRestoreMemory_io_dataRead : 6'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 224:45]
  assign backBufferRestoreMemory_clock = clock;
  assign backBufferRestoreMemory_io_address = backMemoryRestoreCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 216:65]
  assign spriteMemories_0_clock = clock;
  assign spriteMemories_0_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_1_clock = clock;
  assign spriteMemories_1_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_2_clock = clock;
  assign spriteMemories_2_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_3_clock = clock;
  assign spriteMemories_3_io_address = _spriteMemories_3_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_4_clock = clock;
  assign spriteMemories_4_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_5_clock = clock;
  assign spriteMemories_5_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_6_clock = clock;
  assign spriteMemories_6_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_7_clock = clock;
  assign spriteMemories_7_io_address = _spriteMemories_7_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_8_clock = clock;
  assign spriteMemories_8_io_address = _spriteMemories_8_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_9_clock = clock;
  assign spriteMemories_9_io_address = _spriteMemories_9_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_10_clock = clock;
  assign spriteMemories_10_io_address = _spriteMemories_10_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_11_clock = clock;
  assign spriteMemories_11_io_address = _spriteMemories_11_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_12_clock = clock;
  assign spriteMemories_12_io_address = _spriteMemories_12_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_13_clock = clock;
  assign spriteMemories_13_io_address = _spriteMemories_13_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_14_clock = clock;
  assign spriteMemories_14_io_address = _spriteMemories_14_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_15_clock = clock;
  assign spriteMemories_15_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_16_clock = clock;
  assign spriteMemories_16_io_address = _spriteMemories_16_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_17_clock = clock;
  assign spriteMemories_17_io_address = _spriteMemories_17_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_18_clock = clock;
  assign spriteMemories_18_io_address = _spriteMemories_18_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_19_clock = clock;
  assign spriteMemories_19_io_address = _spriteMemories_19_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_20_clock = clock;
  assign spriteMemories_20_io_address = _spriteMemories_20_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_21_clock = clock;
  assign spriteMemories_21_io_address = _spriteMemories_21_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_22_clock = clock;
  assign spriteMemories_22_io_address = _spriteMemories_22_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_23_clock = clock;
  assign spriteMemories_23_io_address = _spriteMemories_23_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_24_clock = clock;
  assign spriteMemories_24_io_address = _spriteMemories_24_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_25_clock = clock;
  assign spriteMemories_25_io_address = _spriteMemories_25_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_26_clock = clock;
  assign spriteMemories_26_io_address = _spriteMemories_26_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_27_clock = clock;
  assign spriteMemories_27_io_address = _spriteMemories_27_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_28_clock = clock;
  assign spriteMemories_28_io_address = _spriteMemories_28_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_29_clock = clock;
  assign spriteMemories_29_io_address = _spriteMemories_29_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_30_clock = clock;
  assign spriteMemories_30_io_address = _spriteMemories_30_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_31_clock = clock;
  assign spriteMemories_31_io_address = _spriteMemories_31_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_32_clock = clock;
  assign spriteMemories_32_io_address = _spriteMemories_32_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_33_clock = clock;
  assign spriteMemories_33_io_address = _spriteMemories_33_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_34_clock = clock;
  assign spriteMemories_34_io_address = _spriteMemories_34_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_35_clock = clock;
  assign spriteMemories_35_io_address = _spriteMemories_35_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_36_clock = clock;
  assign spriteMemories_36_io_address = _spriteMemories_36_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_37_clock = clock;
  assign spriteMemories_37_io_address = _spriteMemories_37_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_38_clock = clock;
  assign spriteMemories_38_io_address = _spriteMemories_38_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_39_clock = clock;
  assign spriteMemories_39_io_address = _spriteMemories_39_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_40_clock = clock;
  assign spriteMemories_40_io_address = _spriteMemories_40_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_41_clock = clock;
  assign spriteMemories_41_io_address = _spriteMemories_41_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_42_clock = clock;
  assign spriteMemories_42_io_address = _spriteMemories_42_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_43_clock = clock;
  assign spriteMemories_43_io_address = _spriteMemories_43_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_44_clock = clock;
  assign spriteMemories_44_io_address = _spriteMemories_44_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_45_clock = clock;
  assign spriteMemories_45_io_address = _spriteMemories_45_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_46_clock = clock;
  assign spriteMemories_46_io_address = _spriteMemories_46_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_47_clock = clock;
  assign spriteMemories_47_io_address = _spriteMemories_47_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_48_clock = clock;
  assign spriteMemories_48_io_address = _spriteMemories_48_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_49_clock = clock;
  assign spriteMemories_49_io_address = _spriteMemories_49_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_50_clock = clock;
  assign spriteMemories_50_io_address = _spriteMemories_50_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_51_clock = clock;
  assign spriteMemories_51_io_address = _spriteMemories_51_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_52_clock = clock;
  assign spriteMemories_52_io_address = _spriteMemories_52_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_53_clock = clock;
  assign spriteMemories_53_io_address = _spriteMemories_53_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_54_clock = clock;
  assign spriteMemories_54_io_address = _spriteMemories_54_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_55_clock = clock;
  assign spriteMemories_55_io_address = _spriteMemories_55_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_56_clock = clock;
  assign spriteMemories_56_io_address = _spriteMemories_56_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_57_clock = clock;
  assign spriteMemories_57_io_address = _spriteMemories_57_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_58_clock = clock;
  assign spriteMemories_58_io_address = _spriteMemories_58_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_59_clock = clock;
  assign spriteMemories_59_io_address = _spriteMemories_59_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_60_clock = clock;
  assign spriteMemories_60_io_address = _spriteMemories_60_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_61_clock = clock;
  assign spriteMemories_61_io_address = _spriteMemories_61_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_62_clock = clock;
  assign spriteMemories_62_io_address = _spriteMemories_62_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_63_clock = clock;
  assign spriteMemories_63_io_address = _spriteMemories_63_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_64_clock = clock;
  assign spriteMemories_64_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_65_clock = clock;
  assign spriteMemories_65_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_66_clock = clock;
  assign spriteMemories_66_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_67_clock = clock;
  assign spriteMemories_67_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_68_clock = clock;
  assign spriteMemories_68_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_69_clock = clock;
  assign spriteMemories_69_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_70_clock = clock;
  assign spriteMemories_70_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_71_clock = clock;
  assign spriteMemories_71_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_72_clock = clock;
  assign spriteMemories_72_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_73_clock = clock;
  assign spriteMemories_73_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_74_clock = clock;
  assign spriteMemories_74_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_75_clock = clock;
  assign spriteMemories_75_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_76_clock = clock;
  assign spriteMemories_76_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_77_clock = clock;
  assign spriteMemories_77_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_78_clock = clock;
  assign spriteMemories_78_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_79_clock = clock;
  assign spriteMemories_79_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_80_clock = clock;
  assign spriteMemories_80_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_81_clock = clock;
  assign spriteMemories_81_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_82_clock = clock;
  assign spriteMemories_82_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_83_clock = clock;
  assign spriteMemories_83_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_84_clock = clock;
  assign spriteMemories_84_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_85_clock = clock;
  assign spriteMemories_85_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_86_clock = clock;
  assign spriteMemories_86_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_87_clock = clock;
  assign spriteMemories_87_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_88_clock = clock;
  assign spriteMemories_88_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_89_clock = clock;
  assign spriteMemories_89_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_90_clock = clock;
  assign spriteMemories_90_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_91_clock = clock;
  assign spriteMemories_91_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_92_clock = clock;
  assign spriteMemories_92_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_93_clock = clock;
  assign spriteMemories_93_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_94_clock = clock;
  assign spriteMemories_94_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_95_clock = clock;
  assign spriteMemories_95_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_96_clock = clock;
  assign spriteMemories_96_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_97_clock = clock;
  assign spriteMemories_97_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_98_clock = clock;
  assign spriteMemories_98_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_99_clock = clock;
  assign spriteMemories_99_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_100_clock = clock;
  assign spriteMemories_100_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_101_clock = clock;
  assign spriteMemories_101_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_102_clock = clock;
  assign spriteMemories_102_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_103_clock = clock;
  assign spriteMemories_103_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_104_clock = clock;
  assign spriteMemories_104_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_105_clock = clock;
  assign spriteMemories_105_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_106_clock = clock;
  assign spriteMemories_106_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_107_clock = clock;
  assign spriteMemories_107_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_108_clock = clock;
  assign spriteMemories_108_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_109_clock = clock;
  assign spriteMemories_109_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_110_clock = clock;
  assign spriteMemories_110_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_111_clock = clock;
  assign spriteMemories_111_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_112_clock = clock;
  assign spriteMemories_112_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_113_clock = clock;
  assign spriteMemories_113_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_114_clock = clock;
  assign spriteMemories_114_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_115_clock = clock;
  assign spriteMemories_115_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_116_clock = clock;
  assign spriteMemories_116_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_117_clock = clock;
  assign spriteMemories_117_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_118_clock = clock;
  assign spriteMemories_118_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_119_clock = clock;
  assign spriteMemories_119_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_120_clock = clock;
  assign spriteMemories_120_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_121_clock = clock;
  assign spriteMemories_121_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_122_clock = clock;
  assign spriteMemories_122_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_123_clock = clock;
  assign spriteMemories_123_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_124_clock = clock;
  assign spriteMemories_124_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_125_clock = clock;
  assign spriteMemories_125_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_126_clock = clock;
  assign spriteMemories_126_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_127_clock = clock;
  assign spriteMemories_127_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign multiHotPriortyReductionTree_io_dataInput_0 = multiHotPriortyReductionTree_io_dataInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_1 = multiHotPriortyReductionTree_io_dataInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_2 = multiHotPriortyReductionTree_io_dataInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_3 = multiHotPriortyReductionTree_io_dataInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_4 = multiHotPriortyReductionTree_io_dataInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_5 = multiHotPriortyReductionTree_io_dataInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_6 = multiHotPriortyReductionTree_io_dataInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_7 = multiHotPriortyReductionTree_io_dataInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_8 = multiHotPriortyReductionTree_io_dataInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_9 = multiHotPriortyReductionTree_io_dataInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_10 = multiHotPriortyReductionTree_io_dataInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_11 = multiHotPriortyReductionTree_io_dataInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_12 = multiHotPriortyReductionTree_io_dataInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_13 = multiHotPriortyReductionTree_io_dataInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_14 = multiHotPriortyReductionTree_io_dataInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_15 = multiHotPriortyReductionTree_io_dataInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_16 = multiHotPriortyReductionTree_io_dataInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_17 = multiHotPriortyReductionTree_io_dataInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_18 = multiHotPriortyReductionTree_io_dataInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_19 = multiHotPriortyReductionTree_io_dataInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_20 = multiHotPriortyReductionTree_io_dataInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_21 = multiHotPriortyReductionTree_io_dataInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_22 = multiHotPriortyReductionTree_io_dataInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_23 = multiHotPriortyReductionTree_io_dataInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_24 = multiHotPriortyReductionTree_io_dataInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_25 = multiHotPriortyReductionTree_io_dataInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_26 = multiHotPriortyReductionTree_io_dataInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_27 = multiHotPriortyReductionTree_io_dataInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_28 = multiHotPriortyReductionTree_io_dataInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_29 = multiHotPriortyReductionTree_io_dataInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_30 = multiHotPriortyReductionTree_io_dataInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_31 = multiHotPriortyReductionTree_io_dataInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_32 = multiHotPriortyReductionTree_io_dataInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_33 = multiHotPriortyReductionTree_io_dataInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_34 = multiHotPriortyReductionTree_io_dataInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_35 = multiHotPriortyReductionTree_io_dataInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_36 = multiHotPriortyReductionTree_io_dataInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_37 = multiHotPriortyReductionTree_io_dataInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_38 = multiHotPriortyReductionTree_io_dataInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_39 = multiHotPriortyReductionTree_io_dataInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_40 = multiHotPriortyReductionTree_io_dataInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_41 = multiHotPriortyReductionTree_io_dataInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_42 = multiHotPriortyReductionTree_io_dataInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_43 = multiHotPriortyReductionTree_io_dataInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_44 = multiHotPriortyReductionTree_io_dataInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_45 = multiHotPriortyReductionTree_io_dataInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_46 = multiHotPriortyReductionTree_io_dataInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_47 = multiHotPriortyReductionTree_io_dataInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_48 = multiHotPriortyReductionTree_io_dataInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_49 = multiHotPriortyReductionTree_io_dataInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_50 = multiHotPriortyReductionTree_io_dataInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_51 = multiHotPriortyReductionTree_io_dataInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_52 = multiHotPriortyReductionTree_io_dataInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_53 = multiHotPriortyReductionTree_io_dataInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_54 = multiHotPriortyReductionTree_io_dataInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_55 = multiHotPriortyReductionTree_io_dataInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_56 = multiHotPriortyReductionTree_io_dataInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_57 = multiHotPriortyReductionTree_io_dataInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_58 = multiHotPriortyReductionTree_io_dataInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_59 = multiHotPriortyReductionTree_io_dataInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_60 = multiHotPriortyReductionTree_io_dataInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_61 = multiHotPriortyReductionTree_io_dataInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_62 = multiHotPriortyReductionTree_io_dataInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_63 = multiHotPriortyReductionTree_io_dataInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_64 = multiHotPriortyReductionTree_io_dataInput_64_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_65 = multiHotPriortyReductionTree_io_dataInput_65_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_66 = multiHotPriortyReductionTree_io_dataInput_66_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_67 = multiHotPriortyReductionTree_io_dataInput_67_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_68 = multiHotPriortyReductionTree_io_dataInput_68_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_69 = multiHotPriortyReductionTree_io_dataInput_69_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_70 = multiHotPriortyReductionTree_io_dataInput_70_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_71 = multiHotPriortyReductionTree_io_dataInput_71_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_72 = multiHotPriortyReductionTree_io_dataInput_72_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_73 = multiHotPriortyReductionTree_io_dataInput_73_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_74 = multiHotPriortyReductionTree_io_dataInput_74_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_75 = multiHotPriortyReductionTree_io_dataInput_75_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_76 = multiHotPriortyReductionTree_io_dataInput_76_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_77 = multiHotPriortyReductionTree_io_dataInput_77_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_78 = multiHotPriortyReductionTree_io_dataInput_78_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_79 = multiHotPriortyReductionTree_io_dataInput_79_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_80 = multiHotPriortyReductionTree_io_dataInput_80_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_81 = multiHotPriortyReductionTree_io_dataInput_81_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_82 = multiHotPriortyReductionTree_io_dataInput_82_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_83 = multiHotPriortyReductionTree_io_dataInput_83_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_84 = multiHotPriortyReductionTree_io_dataInput_84_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_85 = multiHotPriortyReductionTree_io_dataInput_85_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_86 = multiHotPriortyReductionTree_io_dataInput_86_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_87 = multiHotPriortyReductionTree_io_dataInput_87_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_88 = multiHotPriortyReductionTree_io_dataInput_88_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_89 = multiHotPriortyReductionTree_io_dataInput_89_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_90 = multiHotPriortyReductionTree_io_dataInput_90_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_91 = multiHotPriortyReductionTree_io_dataInput_91_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_92 = multiHotPriortyReductionTree_io_dataInput_92_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_93 = multiHotPriortyReductionTree_io_dataInput_93_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_94 = multiHotPriortyReductionTree_io_dataInput_94_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_95 = multiHotPriortyReductionTree_io_dataInput_95_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_96 = multiHotPriortyReductionTree_io_dataInput_96_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_97 = multiHotPriortyReductionTree_io_dataInput_97_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_98 = multiHotPriortyReductionTree_io_dataInput_98_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_99 = multiHotPriortyReductionTree_io_dataInput_99_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_100 = multiHotPriortyReductionTree_io_dataInput_100_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_101 = multiHotPriortyReductionTree_io_dataInput_101_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_102 = multiHotPriortyReductionTree_io_dataInput_102_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_103 = multiHotPriortyReductionTree_io_dataInput_103_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_104 = multiHotPriortyReductionTree_io_dataInput_104_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_105 = multiHotPriortyReductionTree_io_dataInput_105_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_106 = multiHotPriortyReductionTree_io_dataInput_106_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_107 = multiHotPriortyReductionTree_io_dataInput_107_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_108 = multiHotPriortyReductionTree_io_dataInput_108_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_109 = multiHotPriortyReductionTree_io_dataInput_109_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_110 = multiHotPriortyReductionTree_io_dataInput_110_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_111 = multiHotPriortyReductionTree_io_dataInput_111_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_112 = multiHotPriortyReductionTree_io_dataInput_112_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_113 = multiHotPriortyReductionTree_io_dataInput_113_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_114 = multiHotPriortyReductionTree_io_dataInput_114_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_115 = multiHotPriortyReductionTree_io_dataInput_115_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_116 = multiHotPriortyReductionTree_io_dataInput_116_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_117 = multiHotPriortyReductionTree_io_dataInput_117_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_118 = multiHotPriortyReductionTree_io_dataInput_118_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_119 = multiHotPriortyReductionTree_io_dataInput_119_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_120 = multiHotPriortyReductionTree_io_dataInput_120_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_121 = multiHotPriortyReductionTree_io_dataInput_121_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_122 = multiHotPriortyReductionTree_io_dataInput_122_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_123 = multiHotPriortyReductionTree_io_dataInput_123_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_124 = multiHotPriortyReductionTree_io_dataInput_124_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_125 = multiHotPriortyReductionTree_io_dataInput_125_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_126 = multiHotPriortyReductionTree_io_dataInput_126_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_127 = multiHotPriortyReductionTree_io_dataInput_127_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_selectInput_0 = multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_1 = multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_2 = multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_3 = multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_4 = multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_5 = multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_6 = multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_7 = multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_8 = multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_9 = multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_10 = multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_11 = multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_12 = multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_13 = multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_14 = multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_15 = multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_16 = multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_17 = multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_18 = multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_19 = multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_20 = multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_21 = multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_22 = multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_23 = multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_24 = multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_25 = multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_26 = multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_27 = multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_28 = multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_29 = multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_30 = multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_31 = multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_32 = multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_33 = multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_34 = multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_35 = multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_36 = multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_37 = multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_38 = multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_39 = multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_40 = multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_41 = multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_42 = multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_43 = multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_44 = multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_45 = multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_46 = multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_47 = multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_48 = multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_49 = multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_50 = multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_51 = multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_52 = multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_53 = multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_54 = multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_55 = multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_56 = multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_57 = multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_58 = multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_59 = multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_60 = multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_61 = multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_62 = multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_63 = multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_64 = multiHotPriortyReductionTree_io_selectInput_64_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_64_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_64_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_65 = multiHotPriortyReductionTree_io_selectInput_65_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_65_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_65_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_66 = multiHotPriortyReductionTree_io_selectInput_66_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_66_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_66_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_67 = multiHotPriortyReductionTree_io_selectInput_67_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_67_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_67_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_68 = multiHotPriortyReductionTree_io_selectInput_68_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_68_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_68_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_69 = multiHotPriortyReductionTree_io_selectInput_69_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_69_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_69_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_70 = multiHotPriortyReductionTree_io_selectInput_70_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_70_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_70_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_71 = multiHotPriortyReductionTree_io_selectInput_71_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_71_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_71_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_72 = multiHotPriortyReductionTree_io_selectInput_72_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_72_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_72_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_73 = multiHotPriortyReductionTree_io_selectInput_73_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_73_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_73_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_74 = multiHotPriortyReductionTree_io_selectInput_74_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_74_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_74_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_75 = multiHotPriortyReductionTree_io_selectInput_75_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_75_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_75_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_76 = multiHotPriortyReductionTree_io_selectInput_76_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_76_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_76_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_77 = multiHotPriortyReductionTree_io_selectInput_77_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_77_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_77_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_78 = multiHotPriortyReductionTree_io_selectInput_78_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_78_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_78_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_79 = multiHotPriortyReductionTree_io_selectInput_79_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_79_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_79_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_80 = multiHotPriortyReductionTree_io_selectInput_80_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_80_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_80_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_81 = multiHotPriortyReductionTree_io_selectInput_81_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_81_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_81_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_82 = multiHotPriortyReductionTree_io_selectInput_82_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_82_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_82_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_83 = multiHotPriortyReductionTree_io_selectInput_83_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_83_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_83_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_84 = multiHotPriortyReductionTree_io_selectInput_84_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_84_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_84_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_85 = multiHotPriortyReductionTree_io_selectInput_85_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_85_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_85_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_86 = multiHotPriortyReductionTree_io_selectInput_86_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_86_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_86_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_87 = multiHotPriortyReductionTree_io_selectInput_87_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_87_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_87_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_88 = multiHotPriortyReductionTree_io_selectInput_88_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_88_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_88_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_89 = multiHotPriortyReductionTree_io_selectInput_89_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_89_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_89_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_90 = multiHotPriortyReductionTree_io_selectInput_90_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_90_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_90_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_91 = multiHotPriortyReductionTree_io_selectInput_91_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_91_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_91_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_92 = multiHotPriortyReductionTree_io_selectInput_92_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_92_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_92_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_93 = multiHotPriortyReductionTree_io_selectInput_93_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_93_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_93_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_94 = multiHotPriortyReductionTree_io_selectInput_94_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_94_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_94_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_95 = multiHotPriortyReductionTree_io_selectInput_95_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_95_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_95_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_96 = multiHotPriortyReductionTree_io_selectInput_96_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_96_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_96_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_97 = multiHotPriortyReductionTree_io_selectInput_97_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_97_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_97_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_98 = multiHotPriortyReductionTree_io_selectInput_98_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_98_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_98_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_99 = multiHotPriortyReductionTree_io_selectInput_99_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_99_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_99_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_100 = multiHotPriortyReductionTree_io_selectInput_100_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_100_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_100_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_101 = multiHotPriortyReductionTree_io_selectInput_101_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_101_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_101_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_102 = multiHotPriortyReductionTree_io_selectInput_102_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_102_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_102_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_103 = multiHotPriortyReductionTree_io_selectInput_103_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_103_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_103_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_104 = multiHotPriortyReductionTree_io_selectInput_104_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_104_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_104_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_105 = multiHotPriortyReductionTree_io_selectInput_105_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_105_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_105_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_106 = multiHotPriortyReductionTree_io_selectInput_106_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_106_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_106_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_107 = multiHotPriortyReductionTree_io_selectInput_107_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_107_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_107_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_108 = multiHotPriortyReductionTree_io_selectInput_108_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_108_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_108_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_109 = multiHotPriortyReductionTree_io_selectInput_109_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_109_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_109_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_110 = multiHotPriortyReductionTree_io_selectInput_110_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_110_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_110_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_111 = multiHotPriortyReductionTree_io_selectInput_111_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_111_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_111_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_112 = multiHotPriortyReductionTree_io_selectInput_112_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_112_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_112_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_113 = multiHotPriortyReductionTree_io_selectInput_113_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_113_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_113_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_114 = multiHotPriortyReductionTree_io_selectInput_114_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_114_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_114_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_115 = multiHotPriortyReductionTree_io_selectInput_115_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_115_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_115_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_116 = multiHotPriortyReductionTree_io_selectInput_116_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_116_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_116_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_117 = multiHotPriortyReductionTree_io_selectInput_117_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_117_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_117_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_118 = multiHotPriortyReductionTree_io_selectInput_118_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_118_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_118_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_119 = multiHotPriortyReductionTree_io_selectInput_119_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_119_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_119_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_120 = multiHotPriortyReductionTree_io_selectInput_120_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_120_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_120_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_121 = multiHotPriortyReductionTree_io_selectInput_121_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_121_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_121_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_122 = multiHotPriortyReductionTree_io_selectInput_122_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_122_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_122_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_123 = multiHotPriortyReductionTree_io_selectInput_123_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_123_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_123_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_124 = multiHotPriortyReductionTree_io_selectInput_124_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_124_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_124_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_125 = multiHotPriortyReductionTree_io_selectInput_125_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_125_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_125_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_126 = multiHotPriortyReductionTree_io_selectInput_126_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_126_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_126_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_127 = multiHotPriortyReductionTree_io_selectInput_127_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_127_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_127_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
      ScaleCounterReg <= 2'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        ScaleCounterReg <= 2'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 75:23]
      end else begin
        ScaleCounterReg <= _ScaleCounterReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 88:23]
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
      CounterXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        if (CounterXReg == 10'h31f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129]
          CounterXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 77:21]
        end else begin
          CounterXReg <= _CounterXReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 85:21]
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
      CounterYReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        if (CounterXReg == 10'h31f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129]
          CounterYReg <= _GEN_0;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
      backMemoryRestoreCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
    end else if (restoreEnabled) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:70]
      backMemoryRestoreCounter <= _backMemoryRestoreCounter_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 206:30]
    end
    io_Hsync_pipeReg_0 <= io_Hsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_1 <= io_Hsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_2 <= io_Hsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_3 <= ~Hsync; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 94:27]
    io_Vsync_pipeReg_0 <= io_Vsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_1 <= io_Vsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_2 <= io_Vsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_3 <= ~Vsync; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 95:27]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
      frameClockCount <= 21'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
    end else if (frameClockCount == 21'h19a27f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 105:25]
      frameClockCount <= 21'h0;
    end else begin
      frameClockCount <= _frameClockCount_T_2;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_3 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_3 <= io_spriteXPosition_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_7 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_7 <= io_spriteXPosition_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_8 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_8 <= io_spriteXPosition_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_9 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_9 <= io_spriteXPosition_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_10 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_10 <= io_spriteXPosition_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_11 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_11 <= io_spriteXPosition_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_12 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_12 <= io_spriteXPosition_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_13 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_13 <= io_spriteXPosition_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_14 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_14 <= io_spriteXPosition_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_16 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_16 <= io_spriteXPosition_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_17 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_17 <= io_spriteXPosition_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_18 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_18 <= io_spriteXPosition_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_19 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_19 <= io_spriteXPosition_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_20 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_20 <= io_spriteXPosition_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_21 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_21 <= io_spriteXPosition_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_22 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_22 <= io_spriteXPosition_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_23 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_23 <= io_spriteXPosition_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_24 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_24 <= io_spriteXPosition_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_25 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_25 <= io_spriteXPosition_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_26 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_26 <= io_spriteXPosition_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_27 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_27 <= io_spriteXPosition_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_28 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_28 <= io_spriteXPosition_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_29 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_29 <= io_spriteXPosition_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_30 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_30 <= io_spriteXPosition_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_31 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_31 <= io_spriteXPosition_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_32 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_32 <= io_spriteXPosition_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_33 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_33 <= io_spriteXPosition_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_34 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_34 <= io_spriteXPosition_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_35 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_35 <= io_spriteXPosition_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_36 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_36 <= io_spriteXPosition_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_37 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_37 <= io_spriteXPosition_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_38 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_38 <= io_spriteXPosition_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_39 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_39 <= io_spriteXPosition_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_40 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_40 <= io_spriteXPosition_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_41 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_41 <= io_spriteXPosition_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_42 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_42 <= io_spriteXPosition_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_43 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_43 <= io_spriteXPosition_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_44 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_44 <= io_spriteXPosition_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_45 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_45 <= io_spriteXPosition_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_46 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_46 <= io_spriteXPosition_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_47 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_47 <= io_spriteXPosition_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_48 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_48 <= io_spriteXPosition_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_49 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_49 <= io_spriteXPosition_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_50 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_50 <= io_spriteXPosition_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_51 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_51 <= io_spriteXPosition_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_52 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_52 <= io_spriteXPosition_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_53 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_53 <= io_spriteXPosition_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_54 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_54 <= io_spriteXPosition_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_55 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_55 <= io_spriteXPosition_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_56 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_56 <= io_spriteXPosition_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_57 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_57 <= io_spriteXPosition_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_58 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_58 <= io_spriteXPosition_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_59 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_59 <= io_spriteXPosition_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_60 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_60 <= io_spriteXPosition_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_61 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_61 <= io_spriteXPosition_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_62 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_62 <= io_spriteXPosition_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_63 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_63 <= io_spriteXPosition_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_3 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_3 <= io_spriteYPosition_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_7 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_7 <= io_spriteYPosition_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_8 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_8 <= io_spriteYPosition_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_9 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_9 <= io_spriteYPosition_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_10 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_10 <= io_spriteYPosition_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_11 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_11 <= io_spriteYPosition_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_12 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_12 <= io_spriteYPosition_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_13 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_13 <= io_spriteYPosition_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_14 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_14 <= io_spriteYPosition_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_16 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_16 <= io_spriteYPosition_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_17 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_17 <= io_spriteYPosition_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_18 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_18 <= io_spriteYPosition_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_19 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_19 <= io_spriteYPosition_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_20 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_20 <= io_spriteYPosition_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_21 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_21 <= io_spriteYPosition_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_22 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_22 <= io_spriteYPosition_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_23 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_23 <= io_spriteYPosition_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_24 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_24 <= io_spriteYPosition_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_25 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_25 <= io_spriteYPosition_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_26 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_26 <= io_spriteYPosition_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_27 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_27 <= io_spriteYPosition_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_28 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_28 <= io_spriteYPosition_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_29 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_29 <= io_spriteYPosition_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_30 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_30 <= io_spriteYPosition_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_31 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_31 <= io_spriteYPosition_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_32 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_32 <= io_spriteYPosition_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_33 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_33 <= io_spriteYPosition_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_34 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_34 <= io_spriteYPosition_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_35 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_35 <= io_spriteYPosition_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_36 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_36 <= io_spriteYPosition_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_37 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_37 <= io_spriteYPosition_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_38 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_38 <= io_spriteYPosition_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_39 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_39 <= io_spriteYPosition_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_40 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_40 <= io_spriteYPosition_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_41 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_41 <= io_spriteYPosition_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_42 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_42 <= io_spriteYPosition_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_43 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_43 <= io_spriteYPosition_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_44 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_44 <= io_spriteYPosition_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_45 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_45 <= io_spriteYPosition_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_46 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_46 <= io_spriteYPosition_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_47 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_47 <= io_spriteYPosition_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_48 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_48 <= io_spriteYPosition_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_49 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_49 <= io_spriteYPosition_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_50 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_50 <= io_spriteYPosition_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_51 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_51 <= io_spriteYPosition_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_52 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_52 <= io_spriteYPosition_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_53 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_53 <= io_spriteYPosition_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_54 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_54 <= io_spriteYPosition_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_55 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_55 <= io_spriteYPosition_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_56 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_56 <= io_spriteYPosition_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_57 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_57 <= io_spriteYPosition_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_58 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_58 <= io_spriteYPosition_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_59 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_59 <= io_spriteYPosition_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_60 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_60 <= io_spriteYPosition_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_61 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_61 <= io_spriteYPosition_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_62 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_62 <= io_spriteYPosition_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_63 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_63 <= io_spriteYPosition_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    spriteVisibleReg_0 <= reset | _GEN_269; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_1 <= reset | _GEN_270; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_2 <= reset | _GEN_271; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_3 <= reset | _GEN_272; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_4 <= reset | _GEN_273; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_5 <= reset | _GEN_274; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_6 <= reset | _GEN_275; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_7 <= reset | _GEN_276; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_8 <= reset | _GEN_277; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_9 <= reset | _GEN_278; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_10 <= reset | _GEN_279; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_11 <= reset | _GEN_280; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_12 <= reset | _GEN_281; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_13 <= reset | _GEN_282; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_14 <= reset | _GEN_283; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_15 <= reset | _GEN_284; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_16 <= reset | _GEN_285; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_17 <= reset | _GEN_286; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_18 <= reset | _GEN_287; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_19 <= reset | _GEN_288; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_20 <= reset | _GEN_289; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_21 <= reset | _GEN_290; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_22 <= reset | _GEN_291; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_23 <= reset | _GEN_292; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_24 <= reset | _GEN_293; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_25 <= reset | _GEN_294; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_26 <= reset | _GEN_295; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_27 <= reset | _GEN_296; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_28 <= reset | _GEN_297; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_29 <= reset | _GEN_298; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_30 <= reset | _GEN_299; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_31 <= reset | _GEN_300; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_32 <= reset | _GEN_301; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_33 <= reset | _GEN_302; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_34 <= reset | _GEN_303; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_35 <= reset | _GEN_304; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_36 <= reset | _GEN_305; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_37 <= reset | _GEN_306; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_38 <= reset | _GEN_307; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_39 <= reset | _GEN_308; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_40 <= reset | _GEN_309; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_41 <= reset | _GEN_310; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_42 <= reset | _GEN_311; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_43 <= reset | _GEN_312; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_44 <= reset | _GEN_313; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_45 <= reset | _GEN_314; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_46 <= reset | _GEN_315; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_47 <= reset | _GEN_316; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_48 <= reset | _GEN_317; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_49 <= reset | _GEN_318; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_50 <= reset | _GEN_319; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_51 <= reset | _GEN_320; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_52 <= reset | _GEN_321; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_53 <= reset | _GEN_322; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_54 <= reset | _GEN_323; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_55 <= reset | _GEN_324; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_56 <= reset | _GEN_325; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_57 <= reset | _GEN_326; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_58 <= reset | _GEN_327; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_59 <= reset | _GEN_328; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_60 <= reset | _GEN_329; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_61 <= reset | _GEN_330; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_62 <= reset | _GEN_331; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_63 <= reset | _GEN_332; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_64 <= reset | _GEN_333; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_65 <= reset | _GEN_334; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_66 <= reset | _GEN_335; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_67 <= reset | _GEN_336; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_68 <= reset | _GEN_337; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_69 <= reset | _GEN_338; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_70 <= reset | _GEN_339; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_71 <= reset | _GEN_340; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_72 <= reset | _GEN_341; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_73 <= reset | _GEN_342; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_74 <= reset | _GEN_343; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_75 <= reset | _GEN_344; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_76 <= reset | _GEN_345; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_77 <= reset | _GEN_346; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_78 <= reset | _GEN_347; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_79 <= reset | _GEN_348; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_80 <= reset | _GEN_349; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_81 <= reset | _GEN_350; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_82 <= reset | _GEN_351; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_83 <= reset | _GEN_352; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_84 <= reset | _GEN_353; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_85 <= reset | _GEN_354; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_86 <= reset | _GEN_355; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_87 <= reset | _GEN_356; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_88 <= reset | _GEN_357; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_89 <= reset | _GEN_358; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_90 <= reset | _GEN_359; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_91 <= reset | _GEN_360; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_92 <= reset | _GEN_361; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_93 <= reset | _GEN_362; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_94 <= reset | _GEN_363; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_95 <= reset | _GEN_364; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_96 <= reset | _GEN_365; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_97 <= reset | _GEN_366; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_98 <= reset | _GEN_367; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_99 <= reset | _GEN_368; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_100 <= reset | _GEN_369; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_101 <= reset | _GEN_370; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_102 <= reset | _GEN_371; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_103 <= reset | _GEN_372; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_104 <= reset | _GEN_373; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_105 <= reset | _GEN_374; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_106 <= reset | _GEN_375; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_107 <= reset | _GEN_376; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_108 <= reset | _GEN_377; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_109 <= reset | _GEN_378; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_110 <= reset | _GEN_379; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_111 <= reset | _GEN_380; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_112 <= reset | _GEN_381; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_113 <= reset | _GEN_382; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_114 <= reset | _GEN_383; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_115 <= reset | _GEN_384; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_116 <= reset | _GEN_385; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_117 <= reset | _GEN_386; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_118 <= reset | _GEN_387; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_119 <= reset | _GEN_388; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_120 <= reset | _GEN_389; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_121 <= reset | _GEN_390; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_122 <= reset | _GEN_391; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_123 <= reset | _GEN_392; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_124 <= reset | _GEN_393; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_125 <= reset | _GEN_394; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_126 <= reset | _GEN_395; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_127 <= reset | _GEN_396; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_16 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_16 <= io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_17 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_17 <= io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_18 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_18 <= io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_19 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_19 <= io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_20 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_20 <= io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_21 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_21 <= io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_22 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_22 <= io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_23 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_23 <= io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_24 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_24 <= io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_25 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_25 <= io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_26 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_26 <= io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_27 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_27 <= io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_28 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_28 <= io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_29 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_29 <= io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_30 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_30 <= io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_31 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_31 <= io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_32 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_32 <= io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_33 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_33 <= io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_34 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_34 <= io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_35 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_35 <= io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_36 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_36 <= io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_37 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_37 <= io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_38 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_38 <= io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_39 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_39 <= io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_40 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_40 <= io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_41 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_41 <= io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_42 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_42 <= io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_43 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_43 <= io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_44 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_44 <= io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_45 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_45 <= io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_58 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_58 <= io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_59 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_59 <= io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_60 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_60 <= io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_16 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_16 <= io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_17 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_17 <= io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_18 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_18 <= io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_19 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_19 <= io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_20 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_20 <= io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_21 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_21 <= io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_22 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_22 <= io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_23 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_23 <= io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_24 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_24 <= io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_25 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_25 <= io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_26 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_26 <= io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_27 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_27 <= io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_28 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_28 <= io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_29 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_29 <= io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_30 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_30 <= io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_31 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_31 <= io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_32 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_32 <= io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_33 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_33 <= io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_34 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_34 <= io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_35 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_35 <= io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_36 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_36 <= io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_37 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_37 <= io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_38 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_38 <= io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_39 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_39 <= io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_40 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_40 <= io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_41 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_41 <= io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_42 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_42 <= io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_43 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_43 <= io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_44 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_44 <= io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_45 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_45 <= io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_58 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_58 <= io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_59 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_59 <= io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_60 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_60 <= io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
      viewBoxXReg <= io_viewBoxX; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
      viewBoxYReg <= 9'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
      viewBoxYReg <= io_viewBoxY; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
      missingFrameErrorReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
    end else begin
      missingFrameErrorReg <= _GEN_1170;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
      viewBoxOutOfRangeErrorReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
    end else begin
      viewBoxOutOfRangeErrorReg <= _GEN_1167;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
      newFrameStikyReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
    end else if (REG) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:37]
      newFrameStikyReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 152:22]
    end else begin
      newFrameStikyReg <= _GEN_1168;
    end
    REG <= io_frameUpdateDone; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:16]
    backTileMemoryDataRead_0_REG <= backTileMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_1_REG <= backTileMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_2_REG <= backTileMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_3_REG <= backTileMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_4_REG <= backTileMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_5_REG <= backTileMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_6_REG <= backTileMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_7_REG <= backTileMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_8_REG <= backTileMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_9_REG <= backTileMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_10_REG <= backTileMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_11_REG <= backTileMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_12_REG <= backTileMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_13_REG <= backTileMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_14_REG <= backTileMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_15_REG <= backTileMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_16_REG <= backTileMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_17_REG <= backTileMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_18_REG <= backTileMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_19_REG <= backTileMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_20_REG <= backTileMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_21_REG <= backTileMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_22_REG <= backTileMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_23_REG <= backTileMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_24_REG <= backTileMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_25_REG <= backTileMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_26_REG <= backTileMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_27_REG <= backTileMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_28_REG <= backTileMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_29_REG <= backTileMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_30_REG <= backTileMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_31_REG <= backTileMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_32_REG <= backTileMemories_32_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_33_REG <= backTileMemories_33_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_34_REG <= backTileMemories_34_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_35_REG <= backTileMemories_35_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_36_REG <= backTileMemories_36_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_37_REG <= backTileMemories_37_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_38_REG <= backTileMemories_38_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_39_REG <= backTileMemories_39_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_40_REG <= backTileMemories_40_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_41_REG <= backTileMemories_41_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_42_REG <= backTileMemories_42_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_43_REG <= backTileMemories_43_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_44_REG <= backTileMemories_44_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_45_REG <= backTileMemories_45_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_46_REG <= backTileMemories_46_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_47_REG <= backTileMemories_47_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_48_REG <= backTileMemories_48_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_49_REG <= backTileMemories_49_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_50_REG <= backTileMemories_50_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_51_REG <= backTileMemories_51_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_52_REG <= backTileMemories_52_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_53_REG <= backTileMemories_53_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_54_REG <= backTileMemories_54_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_55_REG <= backTileMemories_55_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_56_REG <= backTileMemories_56_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_57_REG <= backTileMemories_57_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_58_REG <= backTileMemories_58_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_59_REG <= backTileMemories_59_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_60_REG <= backTileMemories_60_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_61_REG <= backTileMemories_61_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_62_REG <= backTileMemories_62_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_63_REG <= backTileMemories_63_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
      backMemoryCopyCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
    end else if (preDisplayArea) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23]
      if (backMemoryCopyCounter < 12'h800) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 187:66]
        backMemoryCopyCounter <= _backMemoryCopyCounter_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 188:29]
      end
    end else begin
      backMemoryCopyCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 197:27]
    end
    copyEnabledReg <= preDisplayArea & _T_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23 198:17]
    backBufferShadowMemory_io_address_REG <= backMemoryRestoreCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:92]
    backBufferShadowMemory_io_writeEnable_REG <= backMemoryRestoreCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:33]
    backBufferMemory_io_address_REG <= backMemoryCopyCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:83]
    fullBackgroundColor_REG <= backBufferMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:56]
    if (fullBackgroundColor[6]) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 244:25]
      pixelColorBack <= 6'h0;
    end else begin
      pixelColorBack <= fullBackgroundColor[5:0];
    end
    multiHotPriortyReductionTree_io_dataInput_0_REG <= spriteMemories_0_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1 <= spriteVisibleReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_0_REG <= spriteMemories_0_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_1_REG <= spriteMemories_1_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1 <= spriteVisibleReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_1_REG <= spriteMemories_1_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_2_REG <= spriteMemories_2_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1 <= spriteVisibleReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_2_REG <= spriteMemories_2_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_3_REG <= spriteMemories_3_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1 <= spriteVisibleReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1 <= inSpriteHorizontal_3 & inSpriteVertical_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_3_REG <= spriteMemories_3_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_4_REG <= spriteMemories_4_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1 <= spriteVisibleReg_4; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_4_REG <= spriteMemories_4_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_5_REG <= spriteMemories_5_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1 <= spriteVisibleReg_5; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_5_REG <= spriteMemories_5_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_6_REG <= spriteMemories_6_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1 <= spriteVisibleReg_6; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_6_REG <= spriteMemories_6_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_7_REG <= spriteMemories_7_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1 <= spriteVisibleReg_7; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1 <= inSpriteHorizontal_7 & inSpriteVertical_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_7_REG <= spriteMemories_7_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_8_REG <= spriteMemories_8_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1 <= spriteVisibleReg_8; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1 <= inSpriteHorizontal_8 & inSpriteVertical_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_8_REG <= spriteMemories_8_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_9_REG <= spriteMemories_9_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1 <= spriteVisibleReg_9; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1 <= inSpriteHorizontal_9 & inSpriteVertical_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_9_REG <= spriteMemories_9_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_10_REG <= spriteMemories_10_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1 <= spriteVisibleReg_10; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1 <= inSpriteHorizontal_10 & inSpriteVertical_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_10_REG <= spriteMemories_10_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_11_REG <= spriteMemories_11_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1 <= spriteVisibleReg_11; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1 <= inSpriteHorizontal_11 & inSpriteVertical_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_11_REG <= spriteMemories_11_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_12_REG <= spriteMemories_12_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1 <= spriteVisibleReg_12; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1 <= inSpriteHorizontal_12 & inSpriteVertical_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_12_REG <= spriteMemories_12_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_13_REG <= spriteMemories_13_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1 <= spriteVisibleReg_13; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1 <= inSpriteHorizontal_13 & inSpriteVertical_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_13_REG <= spriteMemories_13_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_14_REG <= spriteMemories_14_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1 <= spriteVisibleReg_14; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1 <= inSpriteHorizontal_14 & inSpriteVertical_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_14_REG <= spriteMemories_14_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_15_REG <= spriteMemories_15_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1 <= spriteVisibleReg_15; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_15_REG <= spriteMemories_15_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_16_REG <= spriteMemories_16_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1 <= spriteVisibleReg_16; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1 <= inSpriteHorizontal_16 & inSpriteVertical_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_16_REG <= spriteMemories_16_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_17_REG <= spriteMemories_17_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1 <= spriteVisibleReg_17; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1 <= inSpriteHorizontal_17 & inSpriteVertical_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_17_REG <= spriteMemories_17_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_18_REG <= spriteMemories_18_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1 <= spriteVisibleReg_18; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1 <= inSpriteHorizontal_18 & inSpriteVertical_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_18_REG <= spriteMemories_18_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_19_REG <= spriteMemories_19_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1 <= spriteVisibleReg_19; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1 <= inSpriteHorizontal_19 & inSpriteVertical_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_19_REG <= spriteMemories_19_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_20_REG <= spriteMemories_20_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1 <= spriteVisibleReg_20; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1 <= inSpriteHorizontal_20 & inSpriteVertical_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_20_REG <= spriteMemories_20_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_21_REG <= spriteMemories_21_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1 <= spriteVisibleReg_21; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1 <= inSpriteHorizontal_21 & inSpriteVertical_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_21_REG <= spriteMemories_21_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_22_REG <= spriteMemories_22_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1 <= spriteVisibleReg_22; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1 <= inSpriteHorizontal_22 & inSpriteVertical_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_22_REG <= spriteMemories_22_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_23_REG <= spriteMemories_23_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1 <= spriteVisibleReg_23; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1 <= inSpriteHorizontal_23 & inSpriteVertical_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_23_REG <= spriteMemories_23_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_24_REG <= spriteMemories_24_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1 <= spriteVisibleReg_24; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1 <= inSpriteHorizontal_24 & inSpriteVertical_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_24_REG <= spriteMemories_24_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_25_REG <= spriteMemories_25_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1 <= spriteVisibleReg_25; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1 <= inSpriteHorizontal_25 & inSpriteVertical_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_25_REG <= spriteMemories_25_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_26_REG <= spriteMemories_26_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1 <= spriteVisibleReg_26; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1 <= inSpriteHorizontal_26 & inSpriteVertical_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_26_REG <= spriteMemories_26_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_27_REG <= spriteMemories_27_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1 <= spriteVisibleReg_27; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1 <= inSpriteHorizontal_27 & inSpriteVertical_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_27_REG <= spriteMemories_27_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_28_REG <= spriteMemories_28_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1 <= spriteVisibleReg_28; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1 <= inSpriteHorizontal_28 & inSpriteVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_28_REG <= spriteMemories_28_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_29_REG <= spriteMemories_29_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1 <= spriteVisibleReg_29; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1 <= inSpriteHorizontal_29 & inSpriteVertical_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_29_REG <= spriteMemories_29_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_30_REG <= spriteMemories_30_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1 <= spriteVisibleReg_30; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1 <= inSpriteHorizontal_30 & inSpriteVertical_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_30_REG <= spriteMemories_30_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_31_REG <= spriteMemories_31_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1 <= spriteVisibleReg_31; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1 <= inSpriteHorizontal_31 & inSpriteVertical_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_31_REG <= spriteMemories_31_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_32_REG <= spriteMemories_32_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1 <= spriteVisibleReg_32; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1 <= inSpriteHorizontal_32 & inSpriteVertical_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_32_REG <= spriteMemories_32_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_33_REG <= spriteMemories_33_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1 <= spriteVisibleReg_33; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1 <= inSpriteHorizontal_33 & inSpriteVertical_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_33_REG <= spriteMemories_33_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_34_REG <= spriteMemories_34_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1 <= spriteVisibleReg_34; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1 <= inSpriteHorizontal_34 & inSpriteVertical_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_34_REG <= spriteMemories_34_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_35_REG <= spriteMemories_35_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1 <= spriteVisibleReg_35; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1 <= inSpriteHorizontal_35 & inSpriteVertical_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_35_REG <= spriteMemories_35_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_36_REG <= spriteMemories_36_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1 <= spriteVisibleReg_36; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1 <= inSpriteHorizontal_36 & inSpriteVertical_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_36_REG <= spriteMemories_36_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_37_REG <= spriteMemories_37_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1 <= spriteVisibleReg_37; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1 <= inSpriteHorizontal_37 & inSpriteVertical_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_37_REG <= spriteMemories_37_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_38_REG <= spriteMemories_38_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1 <= spriteVisibleReg_38; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1 <= inSpriteHorizontal_38 & inSpriteVertical_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_38_REG <= spriteMemories_38_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_39_REG <= spriteMemories_39_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1 <= spriteVisibleReg_39; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1 <= inSpriteHorizontal_39 & inSpriteVertical_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_39_REG <= spriteMemories_39_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_40_REG <= spriteMemories_40_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1 <= spriteVisibleReg_40; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1 <= inSpriteHorizontal_40 & inSpriteVertical_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_40_REG <= spriteMemories_40_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_41_REG <= spriteMemories_41_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1 <= spriteVisibleReg_41; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1 <= inSpriteHorizontal_41 & inSpriteVertical_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_41_REG <= spriteMemories_41_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_42_REG <= spriteMemories_42_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1 <= spriteVisibleReg_42; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1 <= inSpriteHorizontal_42 & inSpriteVertical_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_42_REG <= spriteMemories_42_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_43_REG <= spriteMemories_43_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1 <= spriteVisibleReg_43; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1 <= inSpriteHorizontal_43 & inSpriteVertical_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_43_REG <= spriteMemories_43_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_44_REG <= spriteMemories_44_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1 <= spriteVisibleReg_44; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1 <= inSpriteHorizontal_44 & inSpriteVertical_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_44_REG <= spriteMemories_44_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_45_REG <= spriteMemories_45_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1 <= spriteVisibleReg_45; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1 <= inSpriteHorizontal_45 & inSpriteVertical_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_45_REG <= spriteMemories_45_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_46_REG <= spriteMemories_46_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1 <= spriteVisibleReg_46; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1 <= inSpriteHorizontal_46 & inSpriteVertical_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_46_REG <= spriteMemories_46_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_47_REG <= spriteMemories_47_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1 <= spriteVisibleReg_47; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1 <= inSpriteHorizontal_47 & inSpriteVertical_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_47_REG <= spriteMemories_47_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_48_REG <= spriteMemories_48_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1 <= spriteVisibleReg_48; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1 <= inSpriteHorizontal_48 & inSpriteVertical_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_48_REG <= spriteMemories_48_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_49_REG <= spriteMemories_49_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1 <= spriteVisibleReg_49; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1 <= inSpriteHorizontal_49 & inSpriteVertical_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_49_REG <= spriteMemories_49_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_50_REG <= spriteMemories_50_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1 <= spriteVisibleReg_50; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1 <= inSpriteHorizontal_50 & inSpriteVertical_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_50_REG <= spriteMemories_50_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_51_REG <= spriteMemories_51_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1 <= spriteVisibleReg_51; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1 <= inSpriteHorizontal_51 & inSpriteVertical_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_51_REG <= spriteMemories_51_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_52_REG <= spriteMemories_52_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1 <= spriteVisibleReg_52; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1 <= inSpriteHorizontal_52 & inSpriteVertical_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_52_REG <= spriteMemories_52_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_53_REG <= spriteMemories_53_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1 <= spriteVisibleReg_53; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1 <= inSpriteHorizontal_53 & inSpriteVertical_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_53_REG <= spriteMemories_53_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_54_REG <= spriteMemories_54_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1 <= spriteVisibleReg_54; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1 <= inSpriteHorizontal_54 & inSpriteVertical_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_54_REG <= spriteMemories_54_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_55_REG <= spriteMemories_55_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1 <= spriteVisibleReg_55; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1 <= inSpriteHorizontal_55 & inSpriteVertical_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_55_REG <= spriteMemories_55_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_56_REG <= spriteMemories_56_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1 <= spriteVisibleReg_56; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1 <= inSpriteHorizontal_56 & inSpriteVertical_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_56_REG <= spriteMemories_56_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_57_REG <= spriteMemories_57_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1 <= spriteVisibleReg_57; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1 <= inSpriteHorizontal_57 & inSpriteVertical_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_57_REG <= spriteMemories_57_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_58_REG <= spriteMemories_58_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1 <= spriteVisibleReg_58; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1 <= inSpriteHorizontal_58 & inSpriteVertical_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_58_REG <= spriteMemories_58_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_59_REG <= spriteMemories_59_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1 <= spriteVisibleReg_59; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1 <= inSpriteHorizontal_59 & inSpriteVertical_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_59_REG <= spriteMemories_59_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_60_REG <= spriteMemories_60_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1 <= spriteVisibleReg_60; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1 <= inSpriteHorizontal_60 & inSpriteVertical_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_60_REG <= spriteMemories_60_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_61_REG <= spriteMemories_61_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1 <= spriteVisibleReg_61; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1 <= inSpriteHorizontal_61 & inSpriteVertical_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_61_REG <= spriteMemories_61_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_62_REG <= spriteMemories_62_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1 <= spriteVisibleReg_62; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1 <= inSpriteHorizontal_62 & inSpriteVertical_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_62_REG <= spriteMemories_62_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_63_REG <= spriteMemories_63_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1 <= spriteVisibleReg_63; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1 <= inSpriteHorizontal_63 & inSpriteVertical_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_63_REG <= spriteMemories_63_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_64_REG <= spriteMemories_64_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_64_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_64_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_64_pipeReg__1 <= spriteVisibleReg_64; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_64_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_64_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_64_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_64_REG <= spriteMemories_64_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_65_REG <= spriteMemories_65_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_65_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_65_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_65_pipeReg__1 <= spriteVisibleReg_65; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_65_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_65_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_65_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_65_REG <= spriteMemories_65_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_66_REG <= spriteMemories_66_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_66_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_66_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_66_pipeReg__1 <= spriteVisibleReg_66; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_66_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_66_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_66_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_66_REG <= spriteMemories_66_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_67_REG <= spriteMemories_67_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_67_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_67_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_67_pipeReg__1 <= spriteVisibleReg_67; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_67_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_67_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_67_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_67_REG <= spriteMemories_67_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_68_REG <= spriteMemories_68_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_68_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_68_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_68_pipeReg__1 <= spriteVisibleReg_68; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_68_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_68_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_68_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_68_REG <= spriteMemories_68_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_69_REG <= spriteMemories_69_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_69_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_69_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_69_pipeReg__1 <= spriteVisibleReg_69; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_69_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_69_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_69_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_69_REG <= spriteMemories_69_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_70_REG <= spriteMemories_70_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_70_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_70_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_70_pipeReg__1 <= spriteVisibleReg_70; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_70_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_70_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_70_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_70_REG <= spriteMemories_70_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_71_REG <= spriteMemories_71_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_71_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_71_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_71_pipeReg__1 <= spriteVisibleReg_71; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_71_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_71_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_71_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_71_REG <= spriteMemories_71_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_72_REG <= spriteMemories_72_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_72_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_72_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_72_pipeReg__1 <= spriteVisibleReg_72; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_72_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_72_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_72_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_72_REG <= spriteMemories_72_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_73_REG <= spriteMemories_73_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_73_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_73_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_73_pipeReg__1 <= spriteVisibleReg_73; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_73_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_73_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_73_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_73_REG <= spriteMemories_73_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_74_REG <= spriteMemories_74_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_74_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_74_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_74_pipeReg__1 <= spriteVisibleReg_74; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_74_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_74_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_74_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_74_REG <= spriteMemories_74_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_75_REG <= spriteMemories_75_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_75_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_75_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_75_pipeReg__1 <= spriteVisibleReg_75; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_75_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_75_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_75_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_75_REG <= spriteMemories_75_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_76_REG <= spriteMemories_76_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_76_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_76_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_76_pipeReg__1 <= spriteVisibleReg_76; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_76_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_76_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_76_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_76_REG <= spriteMemories_76_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_77_REG <= spriteMemories_77_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_77_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_77_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_77_pipeReg__1 <= spriteVisibleReg_77; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_77_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_77_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_77_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_77_REG <= spriteMemories_77_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_78_REG <= spriteMemories_78_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_78_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_78_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_78_pipeReg__1 <= spriteVisibleReg_78; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_78_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_78_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_78_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_78_REG <= spriteMemories_78_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_79_REG <= spriteMemories_79_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_79_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_79_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_79_pipeReg__1 <= spriteVisibleReg_79; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_79_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_79_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_79_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_79_REG <= spriteMemories_79_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_80_REG <= spriteMemories_80_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_80_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_80_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_80_pipeReg__1 <= spriteVisibleReg_80; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_80_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_80_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_80_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_80_REG <= spriteMemories_80_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_81_REG <= spriteMemories_81_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_81_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_81_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_81_pipeReg__1 <= spriteVisibleReg_81; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_81_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_81_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_81_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_81_REG <= spriteMemories_81_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_82_REG <= spriteMemories_82_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_82_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_82_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_82_pipeReg__1 <= spriteVisibleReg_82; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_82_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_82_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_82_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_82_REG <= spriteMemories_82_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_83_REG <= spriteMemories_83_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_83_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_83_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_83_pipeReg__1 <= spriteVisibleReg_83; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_83_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_83_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_83_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_83_REG <= spriteMemories_83_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_84_REG <= spriteMemories_84_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_84_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_84_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_84_pipeReg__1 <= spriteVisibleReg_84; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_84_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_84_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_84_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_84_REG <= spriteMemories_84_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_85_REG <= spriteMemories_85_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_85_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_85_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_85_pipeReg__1 <= spriteVisibleReg_85; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_85_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_85_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_85_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_85_REG <= spriteMemories_85_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_86_REG <= spriteMemories_86_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_86_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_86_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_86_pipeReg__1 <= spriteVisibleReg_86; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_86_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_86_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_86_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_86_REG <= spriteMemories_86_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_87_REG <= spriteMemories_87_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_87_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_87_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_87_pipeReg__1 <= spriteVisibleReg_87; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_87_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_87_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_87_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_87_REG <= spriteMemories_87_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_88_REG <= spriteMemories_88_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_88_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_88_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_88_pipeReg__1 <= spriteVisibleReg_88; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_88_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_88_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_88_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_88_REG <= spriteMemories_88_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_89_REG <= spriteMemories_89_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_89_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_89_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_89_pipeReg__1 <= spriteVisibleReg_89; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_89_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_89_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_89_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_89_REG <= spriteMemories_89_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_90_REG <= spriteMemories_90_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_90_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_90_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_90_pipeReg__1 <= spriteVisibleReg_90; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_90_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_90_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_90_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_90_REG <= spriteMemories_90_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_91_REG <= spriteMemories_91_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_91_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_91_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_91_pipeReg__1 <= spriteVisibleReg_91; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_91_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_91_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_91_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_91_REG <= spriteMemories_91_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_92_REG <= spriteMemories_92_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_92_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_92_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_92_pipeReg__1 <= spriteVisibleReg_92; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_92_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_92_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_92_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_92_REG <= spriteMemories_92_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_93_REG <= spriteMemories_93_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_93_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_93_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_93_pipeReg__1 <= spriteVisibleReg_93; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_93_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_93_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_93_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_93_REG <= spriteMemories_93_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_94_REG <= spriteMemories_94_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_94_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_94_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_94_pipeReg__1 <= spriteVisibleReg_94; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_94_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_94_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_94_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_94_REG <= spriteMemories_94_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_95_REG <= spriteMemories_95_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_95_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_95_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_95_pipeReg__1 <= spriteVisibleReg_95; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_95_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_95_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_95_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_95_REG <= spriteMemories_95_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_96_REG <= spriteMemories_96_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_96_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_96_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_96_pipeReg__1 <= spriteVisibleReg_96; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_96_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_96_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_96_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_96_REG <= spriteMemories_96_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_97_REG <= spriteMemories_97_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_97_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_97_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_97_pipeReg__1 <= spriteVisibleReg_97; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_97_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_97_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_97_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_97_REG <= spriteMemories_97_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_98_REG <= spriteMemories_98_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_98_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_98_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_98_pipeReg__1 <= spriteVisibleReg_98; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_98_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_98_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_98_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_98_REG <= spriteMemories_98_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_99_REG <= spriteMemories_99_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_99_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_99_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_99_pipeReg__1 <= spriteVisibleReg_99; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_99_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_99_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_99_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_99_REG <= spriteMemories_99_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_100_REG <= spriteMemories_100_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_100_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_100_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_100_pipeReg__1 <= spriteVisibleReg_100; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_100_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_100_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_100_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_100_REG <= spriteMemories_100_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_101_REG <= spriteMemories_101_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_101_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_101_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_101_pipeReg__1 <= spriteVisibleReg_101; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_101_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_101_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_101_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_101_REG <= spriteMemories_101_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_102_REG <= spriteMemories_102_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_102_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_102_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_102_pipeReg__1 <= spriteVisibleReg_102; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_102_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_102_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_102_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_102_REG <= spriteMemories_102_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_103_REG <= spriteMemories_103_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_103_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_103_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_103_pipeReg__1 <= spriteVisibleReg_103; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_103_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_103_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_103_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_103_REG <= spriteMemories_103_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_104_REG <= spriteMemories_104_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_104_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_104_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_104_pipeReg__1 <= spriteVisibleReg_104; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_104_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_104_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_104_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_104_REG <= spriteMemories_104_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_105_REG <= spriteMemories_105_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_105_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_105_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_105_pipeReg__1 <= spriteVisibleReg_105; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_105_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_105_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_105_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_105_REG <= spriteMemories_105_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_106_REG <= spriteMemories_106_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_106_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_106_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_106_pipeReg__1 <= spriteVisibleReg_106; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_106_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_106_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_106_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_106_REG <= spriteMemories_106_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_107_REG <= spriteMemories_107_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_107_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_107_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_107_pipeReg__1 <= spriteVisibleReg_107; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_107_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_107_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_107_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_107_REG <= spriteMemories_107_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_108_REG <= spriteMemories_108_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_108_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_108_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_108_pipeReg__1 <= spriteVisibleReg_108; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_108_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_108_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_108_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_108_REG <= spriteMemories_108_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_109_REG <= spriteMemories_109_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_109_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_109_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_109_pipeReg__1 <= spriteVisibleReg_109; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_109_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_109_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_109_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_109_REG <= spriteMemories_109_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_110_REG <= spriteMemories_110_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_110_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_110_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_110_pipeReg__1 <= spriteVisibleReg_110; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_110_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_110_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_110_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_110_REG <= spriteMemories_110_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_111_REG <= spriteMemories_111_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_111_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_111_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_111_pipeReg__1 <= spriteVisibleReg_111; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_111_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_111_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_111_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_111_REG <= spriteMemories_111_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_112_REG <= spriteMemories_112_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_112_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_112_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_112_pipeReg__1 <= spriteVisibleReg_112; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_112_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_112_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_112_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_112_REG <= spriteMemories_112_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_113_REG <= spriteMemories_113_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_113_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_113_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_113_pipeReg__1 <= spriteVisibleReg_113; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_113_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_113_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_113_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_113_REG <= spriteMemories_113_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_114_REG <= spriteMemories_114_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_114_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_114_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_114_pipeReg__1 <= spriteVisibleReg_114; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_114_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_114_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_114_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_114_REG <= spriteMemories_114_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_115_REG <= spriteMemories_115_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_115_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_115_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_115_pipeReg__1 <= spriteVisibleReg_115; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_115_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_115_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_115_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_115_REG <= spriteMemories_115_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_116_REG <= spriteMemories_116_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_116_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_116_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_116_pipeReg__1 <= spriteVisibleReg_116; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_116_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_116_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_116_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_116_REG <= spriteMemories_116_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_117_REG <= spriteMemories_117_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_117_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_117_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_117_pipeReg__1 <= spriteVisibleReg_117; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_117_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_117_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_117_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_117_REG <= spriteMemories_117_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_118_REG <= spriteMemories_118_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_118_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_118_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_118_pipeReg__1 <= spriteVisibleReg_118; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_118_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_118_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_118_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_118_REG <= spriteMemories_118_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_119_REG <= spriteMemories_119_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_119_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_119_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_119_pipeReg__1 <= spriteVisibleReg_119; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_119_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_119_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_119_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_119_REG <= spriteMemories_119_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_120_REG <= spriteMemories_120_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_120_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_120_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_120_pipeReg__1 <= spriteVisibleReg_120; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_120_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_120_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_120_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_120_REG <= spriteMemories_120_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_121_REG <= spriteMemories_121_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_121_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_121_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_121_pipeReg__1 <= spriteVisibleReg_121; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_121_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_121_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_121_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_121_REG <= spriteMemories_121_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_122_REG <= spriteMemories_122_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_122_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_122_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_122_pipeReg__1 <= spriteVisibleReg_122; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_122_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_122_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_122_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_122_REG <= spriteMemories_122_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_123_REG <= spriteMemories_123_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_123_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_123_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_123_pipeReg__1 <= spriteVisibleReg_123; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_123_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_123_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_123_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_123_REG <= spriteMemories_123_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_124_REG <= spriteMemories_124_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_124_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_124_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_124_pipeReg__1 <= spriteVisibleReg_124; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_124_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_124_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_124_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_124_REG <= spriteMemories_124_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_125_REG <= spriteMemories_125_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_125_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_125_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_125_pipeReg__1 <= spriteVisibleReg_125; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_125_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_125_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_125_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_125_REG <= spriteMemories_125_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_126_REG <= spriteMemories_126_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_126_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_126_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_126_pipeReg__1 <= spriteVisibleReg_126; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_126_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_126_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_126_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_126_REG <= spriteMemories_126_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_127_REG <= spriteMemories_127_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_127_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_127_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_127_pipeReg__1 <= spriteVisibleReg_127; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_127_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_127_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_127_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_127_REG <= spriteMemories_127_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    pixelColorSprite <= multiHotPriortyReductionTree_io_dataOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 339:33]
    pixelColorSpriteValid <= multiHotPriortyReductionTree_io_selectOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 340:38]
    pixelColourVGA_pipeReg_0 <= pixelColourVGA_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    pixelColourVGA_pipeReg_1 <= pixelColourVGA_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    pixelColourVGA_pipeReg_2 <= CounterXReg < 10'h280 & CounterYReg < 10'h1e0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 97:60]
    io_vgaRed_REG <= {pixelColourVGA[5:4],pixelColourVGA[5:4]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 346:26]
    io_vgaGreen_REG <= {pixelColourVGA[3:2],pixelColourVGA[3:2]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 347:28]
    io_vgaBlue_REG <= {pixelColourVGA[1:0],pixelColourVGA[1:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 348:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ScaleCounterReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  CounterXReg = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  CounterYReg = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  backMemoryRestoreCounter = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  io_Hsync_pipeReg_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_Hsync_pipeReg_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_Hsync_pipeReg_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_Hsync_pipeReg_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_Vsync_pipeReg_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  io_Vsync_pipeReg_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_Vsync_pipeReg_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_Vsync_pipeReg_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  frameClockCount = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXPositionReg_3 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXPositionReg_7 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXPositionReg_8 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXPositionReg_9 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXPositionReg_10 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXPositionReg_11 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXPositionReg_12 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteXPositionReg_13 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  spriteXPositionReg_14 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  spriteXPositionReg_16 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  spriteXPositionReg_17 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  spriteXPositionReg_18 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  spriteXPositionReg_19 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  spriteXPositionReg_20 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  spriteXPositionReg_21 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  spriteXPositionReg_22 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  spriteXPositionReg_23 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  spriteXPositionReg_24 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  spriteXPositionReg_25 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  spriteXPositionReg_26 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  spriteXPositionReg_27 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  spriteXPositionReg_28 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  spriteXPositionReg_29 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  spriteXPositionReg_30 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  spriteXPositionReg_31 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  spriteXPositionReg_32 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  spriteXPositionReg_33 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  spriteXPositionReg_34 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  spriteXPositionReg_35 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  spriteXPositionReg_36 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  spriteXPositionReg_37 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  spriteXPositionReg_38 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  spriteXPositionReg_39 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  spriteXPositionReg_40 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  spriteXPositionReg_41 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  spriteXPositionReg_42 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  spriteXPositionReg_43 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  spriteXPositionReg_44 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  spriteXPositionReg_45 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  spriteXPositionReg_46 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  spriteXPositionReg_47 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  spriteXPositionReg_48 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  spriteXPositionReg_49 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  spriteXPositionReg_50 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  spriteXPositionReg_51 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  spriteXPositionReg_52 = _RAND_58[10:0];
  _RAND_59 = {1{`RANDOM}};
  spriteXPositionReg_53 = _RAND_59[10:0];
  _RAND_60 = {1{`RANDOM}};
  spriteXPositionReg_54 = _RAND_60[10:0];
  _RAND_61 = {1{`RANDOM}};
  spriteXPositionReg_55 = _RAND_61[10:0];
  _RAND_62 = {1{`RANDOM}};
  spriteXPositionReg_56 = _RAND_62[10:0];
  _RAND_63 = {1{`RANDOM}};
  spriteXPositionReg_57 = _RAND_63[10:0];
  _RAND_64 = {1{`RANDOM}};
  spriteXPositionReg_58 = _RAND_64[10:0];
  _RAND_65 = {1{`RANDOM}};
  spriteXPositionReg_59 = _RAND_65[10:0];
  _RAND_66 = {1{`RANDOM}};
  spriteXPositionReg_60 = _RAND_66[10:0];
  _RAND_67 = {1{`RANDOM}};
  spriteXPositionReg_61 = _RAND_67[10:0];
  _RAND_68 = {1{`RANDOM}};
  spriteXPositionReg_62 = _RAND_68[10:0];
  _RAND_69 = {1{`RANDOM}};
  spriteXPositionReg_63 = _RAND_69[10:0];
  _RAND_70 = {1{`RANDOM}};
  spriteYPositionReg_3 = _RAND_70[9:0];
  _RAND_71 = {1{`RANDOM}};
  spriteYPositionReg_7 = _RAND_71[9:0];
  _RAND_72 = {1{`RANDOM}};
  spriteYPositionReg_8 = _RAND_72[9:0];
  _RAND_73 = {1{`RANDOM}};
  spriteYPositionReg_9 = _RAND_73[9:0];
  _RAND_74 = {1{`RANDOM}};
  spriteYPositionReg_10 = _RAND_74[9:0];
  _RAND_75 = {1{`RANDOM}};
  spriteYPositionReg_11 = _RAND_75[9:0];
  _RAND_76 = {1{`RANDOM}};
  spriteYPositionReg_12 = _RAND_76[9:0];
  _RAND_77 = {1{`RANDOM}};
  spriteYPositionReg_13 = _RAND_77[9:0];
  _RAND_78 = {1{`RANDOM}};
  spriteYPositionReg_14 = _RAND_78[9:0];
  _RAND_79 = {1{`RANDOM}};
  spriteYPositionReg_16 = _RAND_79[9:0];
  _RAND_80 = {1{`RANDOM}};
  spriteYPositionReg_17 = _RAND_80[9:0];
  _RAND_81 = {1{`RANDOM}};
  spriteYPositionReg_18 = _RAND_81[9:0];
  _RAND_82 = {1{`RANDOM}};
  spriteYPositionReg_19 = _RAND_82[9:0];
  _RAND_83 = {1{`RANDOM}};
  spriteYPositionReg_20 = _RAND_83[9:0];
  _RAND_84 = {1{`RANDOM}};
  spriteYPositionReg_21 = _RAND_84[9:0];
  _RAND_85 = {1{`RANDOM}};
  spriteYPositionReg_22 = _RAND_85[9:0];
  _RAND_86 = {1{`RANDOM}};
  spriteYPositionReg_23 = _RAND_86[9:0];
  _RAND_87 = {1{`RANDOM}};
  spriteYPositionReg_24 = _RAND_87[9:0];
  _RAND_88 = {1{`RANDOM}};
  spriteYPositionReg_25 = _RAND_88[9:0];
  _RAND_89 = {1{`RANDOM}};
  spriteYPositionReg_26 = _RAND_89[9:0];
  _RAND_90 = {1{`RANDOM}};
  spriteYPositionReg_27 = _RAND_90[9:0];
  _RAND_91 = {1{`RANDOM}};
  spriteYPositionReg_28 = _RAND_91[9:0];
  _RAND_92 = {1{`RANDOM}};
  spriteYPositionReg_29 = _RAND_92[9:0];
  _RAND_93 = {1{`RANDOM}};
  spriteYPositionReg_30 = _RAND_93[9:0];
  _RAND_94 = {1{`RANDOM}};
  spriteYPositionReg_31 = _RAND_94[9:0];
  _RAND_95 = {1{`RANDOM}};
  spriteYPositionReg_32 = _RAND_95[9:0];
  _RAND_96 = {1{`RANDOM}};
  spriteYPositionReg_33 = _RAND_96[9:0];
  _RAND_97 = {1{`RANDOM}};
  spriteYPositionReg_34 = _RAND_97[9:0];
  _RAND_98 = {1{`RANDOM}};
  spriteYPositionReg_35 = _RAND_98[9:0];
  _RAND_99 = {1{`RANDOM}};
  spriteYPositionReg_36 = _RAND_99[9:0];
  _RAND_100 = {1{`RANDOM}};
  spriteYPositionReg_37 = _RAND_100[9:0];
  _RAND_101 = {1{`RANDOM}};
  spriteYPositionReg_38 = _RAND_101[9:0];
  _RAND_102 = {1{`RANDOM}};
  spriteYPositionReg_39 = _RAND_102[9:0];
  _RAND_103 = {1{`RANDOM}};
  spriteYPositionReg_40 = _RAND_103[9:0];
  _RAND_104 = {1{`RANDOM}};
  spriteYPositionReg_41 = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  spriteYPositionReg_42 = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  spriteYPositionReg_43 = _RAND_106[9:0];
  _RAND_107 = {1{`RANDOM}};
  spriteYPositionReg_44 = _RAND_107[9:0];
  _RAND_108 = {1{`RANDOM}};
  spriteYPositionReg_45 = _RAND_108[9:0];
  _RAND_109 = {1{`RANDOM}};
  spriteYPositionReg_46 = _RAND_109[9:0];
  _RAND_110 = {1{`RANDOM}};
  spriteYPositionReg_47 = _RAND_110[9:0];
  _RAND_111 = {1{`RANDOM}};
  spriteYPositionReg_48 = _RAND_111[9:0];
  _RAND_112 = {1{`RANDOM}};
  spriteYPositionReg_49 = _RAND_112[9:0];
  _RAND_113 = {1{`RANDOM}};
  spriteYPositionReg_50 = _RAND_113[9:0];
  _RAND_114 = {1{`RANDOM}};
  spriteYPositionReg_51 = _RAND_114[9:0];
  _RAND_115 = {1{`RANDOM}};
  spriteYPositionReg_52 = _RAND_115[9:0];
  _RAND_116 = {1{`RANDOM}};
  spriteYPositionReg_53 = _RAND_116[9:0];
  _RAND_117 = {1{`RANDOM}};
  spriteYPositionReg_54 = _RAND_117[9:0];
  _RAND_118 = {1{`RANDOM}};
  spriteYPositionReg_55 = _RAND_118[9:0];
  _RAND_119 = {1{`RANDOM}};
  spriteYPositionReg_56 = _RAND_119[9:0];
  _RAND_120 = {1{`RANDOM}};
  spriteYPositionReg_57 = _RAND_120[9:0];
  _RAND_121 = {1{`RANDOM}};
  spriteYPositionReg_58 = _RAND_121[9:0];
  _RAND_122 = {1{`RANDOM}};
  spriteYPositionReg_59 = _RAND_122[9:0];
  _RAND_123 = {1{`RANDOM}};
  spriteYPositionReg_60 = _RAND_123[9:0];
  _RAND_124 = {1{`RANDOM}};
  spriteYPositionReg_61 = _RAND_124[9:0];
  _RAND_125 = {1{`RANDOM}};
  spriteYPositionReg_62 = _RAND_125[9:0];
  _RAND_126 = {1{`RANDOM}};
  spriteYPositionReg_63 = _RAND_126[9:0];
  _RAND_127 = {1{`RANDOM}};
  spriteVisibleReg_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  spriteVisibleReg_1 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  spriteVisibleReg_2 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  spriteVisibleReg_3 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  spriteVisibleReg_4 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  spriteVisibleReg_5 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  spriteVisibleReg_6 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  spriteVisibleReg_7 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  spriteVisibleReg_8 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  spriteVisibleReg_9 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  spriteVisibleReg_10 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  spriteVisibleReg_11 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  spriteVisibleReg_12 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  spriteVisibleReg_13 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  spriteVisibleReg_14 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  spriteVisibleReg_15 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  spriteVisibleReg_16 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  spriteVisibleReg_17 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  spriteVisibleReg_18 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  spriteVisibleReg_19 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  spriteVisibleReg_20 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  spriteVisibleReg_21 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  spriteVisibleReg_22 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  spriteVisibleReg_23 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  spriteVisibleReg_24 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  spriteVisibleReg_25 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  spriteVisibleReg_26 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  spriteVisibleReg_27 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  spriteVisibleReg_28 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  spriteVisibleReg_29 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  spriteVisibleReg_30 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  spriteVisibleReg_31 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  spriteVisibleReg_32 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  spriteVisibleReg_33 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  spriteVisibleReg_34 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  spriteVisibleReg_35 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  spriteVisibleReg_36 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  spriteVisibleReg_37 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  spriteVisibleReg_38 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  spriteVisibleReg_39 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  spriteVisibleReg_40 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  spriteVisibleReg_41 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  spriteVisibleReg_42 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  spriteVisibleReg_43 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  spriteVisibleReg_44 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  spriteVisibleReg_45 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  spriteVisibleReg_46 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  spriteVisibleReg_47 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  spriteVisibleReg_48 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  spriteVisibleReg_49 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  spriteVisibleReg_50 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  spriteVisibleReg_51 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  spriteVisibleReg_52 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  spriteVisibleReg_53 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  spriteVisibleReg_54 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  spriteVisibleReg_55 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  spriteVisibleReg_56 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  spriteVisibleReg_57 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  spriteVisibleReg_58 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  spriteVisibleReg_59 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  spriteVisibleReg_60 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  spriteVisibleReg_61 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  spriteVisibleReg_62 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  spriteVisibleReg_63 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  spriteVisibleReg_64 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  spriteVisibleReg_65 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  spriteVisibleReg_66 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  spriteVisibleReg_67 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  spriteVisibleReg_68 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  spriteVisibleReg_69 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  spriteVisibleReg_70 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  spriteVisibleReg_71 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  spriteVisibleReg_72 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  spriteVisibleReg_73 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  spriteVisibleReg_74 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  spriteVisibleReg_75 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  spriteVisibleReg_76 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  spriteVisibleReg_77 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  spriteVisibleReg_78 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  spriteVisibleReg_79 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  spriteVisibleReg_80 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  spriteVisibleReg_81 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  spriteVisibleReg_82 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  spriteVisibleReg_83 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  spriteVisibleReg_84 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  spriteVisibleReg_85 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  spriteVisibleReg_86 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  spriteVisibleReg_87 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  spriteVisibleReg_88 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  spriteVisibleReg_89 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  spriteVisibleReg_90 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  spriteVisibleReg_91 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  spriteVisibleReg_92 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  spriteVisibleReg_93 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  spriteVisibleReg_94 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  spriteVisibleReg_95 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  spriteVisibleReg_96 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  spriteVisibleReg_97 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  spriteVisibleReg_98 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  spriteVisibleReg_99 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  spriteVisibleReg_100 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  spriteVisibleReg_101 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  spriteVisibleReg_102 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  spriteVisibleReg_103 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  spriteVisibleReg_104 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  spriteVisibleReg_105 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  spriteVisibleReg_106 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  spriteVisibleReg_107 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  spriteVisibleReg_108 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  spriteVisibleReg_109 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  spriteVisibleReg_110 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  spriteVisibleReg_111 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  spriteVisibleReg_112 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  spriteVisibleReg_113 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  spriteVisibleReg_114 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  spriteVisibleReg_115 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  spriteVisibleReg_116 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  spriteVisibleReg_117 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  spriteVisibleReg_118 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  spriteVisibleReg_119 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  spriteVisibleReg_120 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  spriteVisibleReg_121 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  spriteVisibleReg_122 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  spriteVisibleReg_123 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  spriteVisibleReg_124 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  spriteVisibleReg_125 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  spriteVisibleReg_126 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  spriteVisibleReg_127 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_16 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_17 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_18 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_19 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_20 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_21 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_22 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_23 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_24 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_25 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_26 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_27 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_28 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_29 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_30 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_31 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_32 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_33 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_34 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_35 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_36 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_37 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_38 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_39 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_40 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_41 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_42 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_43 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_44 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_45 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_58 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_59 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_60 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_16 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_17 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_18 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_19 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_20 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_21 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_22 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_23 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_24 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_25 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_26 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_27 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_28 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_29 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_30 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_31 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_32 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_33 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_34 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_35 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_36 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_37 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_38 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_39 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_40 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_41 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_42 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_43 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_44 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_45 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_58 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_59 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_60 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  viewBoxXReg = _RAND_321[9:0];
  _RAND_322 = {1{`RANDOM}};
  viewBoxYReg = _RAND_322[8:0];
  _RAND_323 = {1{`RANDOM}};
  missingFrameErrorReg = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  viewBoxOutOfRangeErrorReg = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  newFrameStikyReg = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  REG = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  backTileMemoryDataRead_0_REG = _RAND_327[6:0];
  _RAND_328 = {1{`RANDOM}};
  backTileMemoryDataRead_1_REG = _RAND_328[6:0];
  _RAND_329 = {1{`RANDOM}};
  backTileMemoryDataRead_2_REG = _RAND_329[6:0];
  _RAND_330 = {1{`RANDOM}};
  backTileMemoryDataRead_3_REG = _RAND_330[6:0];
  _RAND_331 = {1{`RANDOM}};
  backTileMemoryDataRead_4_REG = _RAND_331[6:0];
  _RAND_332 = {1{`RANDOM}};
  backTileMemoryDataRead_5_REG = _RAND_332[6:0];
  _RAND_333 = {1{`RANDOM}};
  backTileMemoryDataRead_6_REG = _RAND_333[6:0];
  _RAND_334 = {1{`RANDOM}};
  backTileMemoryDataRead_7_REG = _RAND_334[6:0];
  _RAND_335 = {1{`RANDOM}};
  backTileMemoryDataRead_8_REG = _RAND_335[6:0];
  _RAND_336 = {1{`RANDOM}};
  backTileMemoryDataRead_9_REG = _RAND_336[6:0];
  _RAND_337 = {1{`RANDOM}};
  backTileMemoryDataRead_10_REG = _RAND_337[6:0];
  _RAND_338 = {1{`RANDOM}};
  backTileMemoryDataRead_11_REG = _RAND_338[6:0];
  _RAND_339 = {1{`RANDOM}};
  backTileMemoryDataRead_12_REG = _RAND_339[6:0];
  _RAND_340 = {1{`RANDOM}};
  backTileMemoryDataRead_13_REG = _RAND_340[6:0];
  _RAND_341 = {1{`RANDOM}};
  backTileMemoryDataRead_14_REG = _RAND_341[6:0];
  _RAND_342 = {1{`RANDOM}};
  backTileMemoryDataRead_15_REG = _RAND_342[6:0];
  _RAND_343 = {1{`RANDOM}};
  backTileMemoryDataRead_16_REG = _RAND_343[6:0];
  _RAND_344 = {1{`RANDOM}};
  backTileMemoryDataRead_17_REG = _RAND_344[6:0];
  _RAND_345 = {1{`RANDOM}};
  backTileMemoryDataRead_18_REG = _RAND_345[6:0];
  _RAND_346 = {1{`RANDOM}};
  backTileMemoryDataRead_19_REG = _RAND_346[6:0];
  _RAND_347 = {1{`RANDOM}};
  backTileMemoryDataRead_20_REG = _RAND_347[6:0];
  _RAND_348 = {1{`RANDOM}};
  backTileMemoryDataRead_21_REG = _RAND_348[6:0];
  _RAND_349 = {1{`RANDOM}};
  backTileMemoryDataRead_22_REG = _RAND_349[6:0];
  _RAND_350 = {1{`RANDOM}};
  backTileMemoryDataRead_23_REG = _RAND_350[6:0];
  _RAND_351 = {1{`RANDOM}};
  backTileMemoryDataRead_24_REG = _RAND_351[6:0];
  _RAND_352 = {1{`RANDOM}};
  backTileMemoryDataRead_25_REG = _RAND_352[6:0];
  _RAND_353 = {1{`RANDOM}};
  backTileMemoryDataRead_26_REG = _RAND_353[6:0];
  _RAND_354 = {1{`RANDOM}};
  backTileMemoryDataRead_27_REG = _RAND_354[6:0];
  _RAND_355 = {1{`RANDOM}};
  backTileMemoryDataRead_28_REG = _RAND_355[6:0];
  _RAND_356 = {1{`RANDOM}};
  backTileMemoryDataRead_29_REG = _RAND_356[6:0];
  _RAND_357 = {1{`RANDOM}};
  backTileMemoryDataRead_30_REG = _RAND_357[6:0];
  _RAND_358 = {1{`RANDOM}};
  backTileMemoryDataRead_31_REG = _RAND_358[6:0];
  _RAND_359 = {1{`RANDOM}};
  backTileMemoryDataRead_32_REG = _RAND_359[6:0];
  _RAND_360 = {1{`RANDOM}};
  backTileMemoryDataRead_33_REG = _RAND_360[6:0];
  _RAND_361 = {1{`RANDOM}};
  backTileMemoryDataRead_34_REG = _RAND_361[6:0];
  _RAND_362 = {1{`RANDOM}};
  backTileMemoryDataRead_35_REG = _RAND_362[6:0];
  _RAND_363 = {1{`RANDOM}};
  backTileMemoryDataRead_36_REG = _RAND_363[6:0];
  _RAND_364 = {1{`RANDOM}};
  backTileMemoryDataRead_37_REG = _RAND_364[6:0];
  _RAND_365 = {1{`RANDOM}};
  backTileMemoryDataRead_38_REG = _RAND_365[6:0];
  _RAND_366 = {1{`RANDOM}};
  backTileMemoryDataRead_39_REG = _RAND_366[6:0];
  _RAND_367 = {1{`RANDOM}};
  backTileMemoryDataRead_40_REG = _RAND_367[6:0];
  _RAND_368 = {1{`RANDOM}};
  backTileMemoryDataRead_41_REG = _RAND_368[6:0];
  _RAND_369 = {1{`RANDOM}};
  backTileMemoryDataRead_42_REG = _RAND_369[6:0];
  _RAND_370 = {1{`RANDOM}};
  backTileMemoryDataRead_43_REG = _RAND_370[6:0];
  _RAND_371 = {1{`RANDOM}};
  backTileMemoryDataRead_44_REG = _RAND_371[6:0];
  _RAND_372 = {1{`RANDOM}};
  backTileMemoryDataRead_45_REG = _RAND_372[6:0];
  _RAND_373 = {1{`RANDOM}};
  backTileMemoryDataRead_46_REG = _RAND_373[6:0];
  _RAND_374 = {1{`RANDOM}};
  backTileMemoryDataRead_47_REG = _RAND_374[6:0];
  _RAND_375 = {1{`RANDOM}};
  backTileMemoryDataRead_48_REG = _RAND_375[6:0];
  _RAND_376 = {1{`RANDOM}};
  backTileMemoryDataRead_49_REG = _RAND_376[6:0];
  _RAND_377 = {1{`RANDOM}};
  backTileMemoryDataRead_50_REG = _RAND_377[6:0];
  _RAND_378 = {1{`RANDOM}};
  backTileMemoryDataRead_51_REG = _RAND_378[6:0];
  _RAND_379 = {1{`RANDOM}};
  backTileMemoryDataRead_52_REG = _RAND_379[6:0];
  _RAND_380 = {1{`RANDOM}};
  backTileMemoryDataRead_53_REG = _RAND_380[6:0];
  _RAND_381 = {1{`RANDOM}};
  backTileMemoryDataRead_54_REG = _RAND_381[6:0];
  _RAND_382 = {1{`RANDOM}};
  backTileMemoryDataRead_55_REG = _RAND_382[6:0];
  _RAND_383 = {1{`RANDOM}};
  backTileMemoryDataRead_56_REG = _RAND_383[6:0];
  _RAND_384 = {1{`RANDOM}};
  backTileMemoryDataRead_57_REG = _RAND_384[6:0];
  _RAND_385 = {1{`RANDOM}};
  backTileMemoryDataRead_58_REG = _RAND_385[6:0];
  _RAND_386 = {1{`RANDOM}};
  backTileMemoryDataRead_59_REG = _RAND_386[6:0];
  _RAND_387 = {1{`RANDOM}};
  backTileMemoryDataRead_60_REG = _RAND_387[6:0];
  _RAND_388 = {1{`RANDOM}};
  backTileMemoryDataRead_61_REG = _RAND_388[6:0];
  _RAND_389 = {1{`RANDOM}};
  backTileMemoryDataRead_62_REG = _RAND_389[6:0];
  _RAND_390 = {1{`RANDOM}};
  backTileMemoryDataRead_63_REG = _RAND_390[6:0];
  _RAND_391 = {1{`RANDOM}};
  backMemoryCopyCounter = _RAND_391[11:0];
  _RAND_392 = {1{`RANDOM}};
  copyEnabledReg = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  backBufferShadowMemory_io_address_REG = _RAND_393[10:0];
  _RAND_394 = {1{`RANDOM}};
  backBufferShadowMemory_io_writeEnable_REG = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  backBufferMemory_io_address_REG = _RAND_395[10:0];
  _RAND_396 = {1{`RANDOM}};
  fullBackgroundColor_REG = _RAND_396[5:0];
  _RAND_397 = {1{`RANDOM}};
  pixelColorBack = _RAND_397[5:0];
  _RAND_398 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_0_REG = _RAND_398[5:0];
  _RAND_399 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_REG = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_1_REG = _RAND_404[5:0];
  _RAND_405 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_REG = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_2_REG = _RAND_410[5:0];
  _RAND_411 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_REG = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_3_REG = _RAND_416[5:0];
  _RAND_417 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_REG = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_4_REG = _RAND_422[5:0];
  _RAND_423 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_REG = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_5_REG = _RAND_428[5:0];
  _RAND_429 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_REG = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_6_REG = _RAND_434[5:0];
  _RAND_435 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_REG = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_7_REG = _RAND_440[5:0];
  _RAND_441 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_REG = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_8_REG = _RAND_446[5:0];
  _RAND_447 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_REG = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_9_REG = _RAND_452[5:0];
  _RAND_453 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_REG = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_10_REG = _RAND_458[5:0];
  _RAND_459 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_REG = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_11_REG = _RAND_464[5:0];
  _RAND_465 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_REG = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_12_REG = _RAND_470[5:0];
  _RAND_471 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_REG = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_13_REG = _RAND_476[5:0];
  _RAND_477 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_REG = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_14_REG = _RAND_482[5:0];
  _RAND_483 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_REG = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_15_REG = _RAND_488[5:0];
  _RAND_489 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_REG = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_16_REG = _RAND_494[5:0];
  _RAND_495 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_REG = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_17_REG = _RAND_500[5:0];
  _RAND_501 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_REG = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_18_REG = _RAND_506[5:0];
  _RAND_507 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_REG = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_19_REG = _RAND_512[5:0];
  _RAND_513 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_REG = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_20_REG = _RAND_518[5:0];
  _RAND_519 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_REG = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_21_REG = _RAND_524[5:0];
  _RAND_525 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_REG = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_22_REG = _RAND_530[5:0];
  _RAND_531 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_REG = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_23_REG = _RAND_536[5:0];
  _RAND_537 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_REG = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_24_REG = _RAND_542[5:0];
  _RAND_543 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_REG = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_25_REG = _RAND_548[5:0];
  _RAND_549 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_REG = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_26_REG = _RAND_554[5:0];
  _RAND_555 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_REG = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_27_REG = _RAND_560[5:0];
  _RAND_561 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_REG = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_28_REG = _RAND_566[5:0];
  _RAND_567 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_REG = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_29_REG = _RAND_572[5:0];
  _RAND_573 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_REG = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_30_REG = _RAND_578[5:0];
  _RAND_579 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_REG = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_31_REG = _RAND_584[5:0];
  _RAND_585 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_REG = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_32_REG = _RAND_590[5:0];
  _RAND_591 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_REG = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_33_REG = _RAND_596[5:0];
  _RAND_597 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_REG = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_34_REG = _RAND_602[5:0];
  _RAND_603 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_REG = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_35_REG = _RAND_608[5:0];
  _RAND_609 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_REG = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_36_REG = _RAND_614[5:0];
  _RAND_615 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_REG = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_37_REG = _RAND_620[5:0];
  _RAND_621 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_REG = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_38_REG = _RAND_626[5:0];
  _RAND_627 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_REG = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_39_REG = _RAND_632[5:0];
  _RAND_633 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_REG = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_40_REG = _RAND_638[5:0];
  _RAND_639 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_REG = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_41_REG = _RAND_644[5:0];
  _RAND_645 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_REG = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_42_REG = _RAND_650[5:0];
  _RAND_651 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_REG = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_43_REG = _RAND_656[5:0];
  _RAND_657 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_REG = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_44_REG = _RAND_662[5:0];
  _RAND_663 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_REG = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_45_REG = _RAND_668[5:0];
  _RAND_669 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_REG = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_46_REG = _RAND_674[5:0];
  _RAND_675 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_REG = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_47_REG = _RAND_680[5:0];
  _RAND_681 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_REG = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_48_REG = _RAND_686[5:0];
  _RAND_687 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_REG = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_49_REG = _RAND_692[5:0];
  _RAND_693 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_REG = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_50_REG = _RAND_698[5:0];
  _RAND_699 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_REG = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_51_REG = _RAND_704[5:0];
  _RAND_705 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_REG = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_52_REG = _RAND_710[5:0];
  _RAND_711 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_REG = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_53_REG = _RAND_716[5:0];
  _RAND_717 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_REG = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_54_REG = _RAND_722[5:0];
  _RAND_723 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_REG = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_55_REG = _RAND_728[5:0];
  _RAND_729 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_REG = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_56_REG = _RAND_734[5:0];
  _RAND_735 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_REG = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_57_REG = _RAND_740[5:0];
  _RAND_741 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_REG = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_58_REG = _RAND_746[5:0];
  _RAND_747 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_REG = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_59_REG = _RAND_752[5:0];
  _RAND_753 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_REG = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_60_REG = _RAND_758[5:0];
  _RAND_759 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_REG = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_61_REG = _RAND_764[5:0];
  _RAND_765 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_REG = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_62_REG = _RAND_770[5:0];
  _RAND_771 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_REG = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_63_REG = _RAND_776[5:0];
  _RAND_777 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_REG = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_64_REG = _RAND_782[5:0];
  _RAND_783 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_64_pipeReg__0 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_64_pipeReg__1 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_64_pipeReg_1_0 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_64_pipeReg_1_1 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_64_REG = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_65_REG = _RAND_788[5:0];
  _RAND_789 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_65_pipeReg__0 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_65_pipeReg__1 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_65_pipeReg_1_0 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_65_pipeReg_1_1 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_65_REG = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_66_REG = _RAND_794[5:0];
  _RAND_795 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_66_pipeReg__0 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_66_pipeReg__1 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_66_pipeReg_1_0 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_66_pipeReg_1_1 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_66_REG = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_67_REG = _RAND_800[5:0];
  _RAND_801 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_67_pipeReg__0 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_67_pipeReg__1 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_67_pipeReg_1_0 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_67_pipeReg_1_1 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_67_REG = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_68_REG = _RAND_806[5:0];
  _RAND_807 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_68_pipeReg__0 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_68_pipeReg__1 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_68_pipeReg_1_0 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_68_pipeReg_1_1 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_68_REG = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_69_REG = _RAND_812[5:0];
  _RAND_813 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_69_pipeReg__0 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_69_pipeReg__1 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_69_pipeReg_1_0 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_69_pipeReg_1_1 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_69_REG = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_70_REG = _RAND_818[5:0];
  _RAND_819 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_70_pipeReg__0 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_70_pipeReg__1 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_70_pipeReg_1_0 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_70_pipeReg_1_1 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_70_REG = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_71_REG = _RAND_824[5:0];
  _RAND_825 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_71_pipeReg__0 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_71_pipeReg__1 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_71_pipeReg_1_0 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_71_pipeReg_1_1 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_71_REG = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_72_REG = _RAND_830[5:0];
  _RAND_831 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_72_pipeReg__0 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_72_pipeReg__1 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_72_pipeReg_1_0 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_72_pipeReg_1_1 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_72_REG = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_73_REG = _RAND_836[5:0];
  _RAND_837 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_73_pipeReg__0 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_73_pipeReg__1 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_73_pipeReg_1_0 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_73_pipeReg_1_1 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_73_REG = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_74_REG = _RAND_842[5:0];
  _RAND_843 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_74_pipeReg__0 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_74_pipeReg__1 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_74_pipeReg_1_0 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_74_pipeReg_1_1 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_74_REG = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_75_REG = _RAND_848[5:0];
  _RAND_849 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_75_pipeReg__0 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_75_pipeReg__1 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_75_pipeReg_1_0 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_75_pipeReg_1_1 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_75_REG = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_76_REG = _RAND_854[5:0];
  _RAND_855 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_76_pipeReg__0 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_76_pipeReg__1 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_76_pipeReg_1_0 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_76_pipeReg_1_1 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_76_REG = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_77_REG = _RAND_860[5:0];
  _RAND_861 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_77_pipeReg__0 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_77_pipeReg__1 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_77_pipeReg_1_0 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_77_pipeReg_1_1 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_77_REG = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_78_REG = _RAND_866[5:0];
  _RAND_867 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_78_pipeReg__0 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_78_pipeReg__1 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_78_pipeReg_1_0 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_78_pipeReg_1_1 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_78_REG = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_79_REG = _RAND_872[5:0];
  _RAND_873 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_79_pipeReg__0 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_79_pipeReg__1 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_79_pipeReg_1_0 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_79_pipeReg_1_1 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_79_REG = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_80_REG = _RAND_878[5:0];
  _RAND_879 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_80_pipeReg__0 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_80_pipeReg__1 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_80_pipeReg_1_0 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_80_pipeReg_1_1 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_80_REG = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_81_REG = _RAND_884[5:0];
  _RAND_885 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_81_pipeReg__0 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_81_pipeReg__1 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_81_pipeReg_1_0 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_81_pipeReg_1_1 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_81_REG = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_82_REG = _RAND_890[5:0];
  _RAND_891 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_82_pipeReg__0 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_82_pipeReg__1 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_82_pipeReg_1_0 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_82_pipeReg_1_1 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_82_REG = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_83_REG = _RAND_896[5:0];
  _RAND_897 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_83_pipeReg__0 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_83_pipeReg__1 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_83_pipeReg_1_0 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_83_pipeReg_1_1 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_83_REG = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_84_REG = _RAND_902[5:0];
  _RAND_903 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_84_pipeReg__0 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_84_pipeReg__1 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_84_pipeReg_1_0 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_84_pipeReg_1_1 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_84_REG = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_85_REG = _RAND_908[5:0];
  _RAND_909 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_85_pipeReg__0 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_85_pipeReg__1 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_85_pipeReg_1_0 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_85_pipeReg_1_1 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_85_REG = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_86_REG = _RAND_914[5:0];
  _RAND_915 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_86_pipeReg__0 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_86_pipeReg__1 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_86_pipeReg_1_0 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_86_pipeReg_1_1 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_86_REG = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_87_REG = _RAND_920[5:0];
  _RAND_921 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_87_pipeReg__0 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_87_pipeReg__1 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_87_pipeReg_1_0 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_87_pipeReg_1_1 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_87_REG = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_88_REG = _RAND_926[5:0];
  _RAND_927 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_88_pipeReg__0 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_88_pipeReg__1 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_88_pipeReg_1_0 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_88_pipeReg_1_1 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_88_REG = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_89_REG = _RAND_932[5:0];
  _RAND_933 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_89_pipeReg__0 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_89_pipeReg__1 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_89_pipeReg_1_0 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_89_pipeReg_1_1 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_89_REG = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_90_REG = _RAND_938[5:0];
  _RAND_939 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_90_pipeReg__0 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_90_pipeReg__1 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_90_pipeReg_1_0 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_90_pipeReg_1_1 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_90_REG = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_91_REG = _RAND_944[5:0];
  _RAND_945 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_91_pipeReg__0 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_91_pipeReg__1 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_91_pipeReg_1_0 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_91_pipeReg_1_1 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_91_REG = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_92_REG = _RAND_950[5:0];
  _RAND_951 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_92_pipeReg__0 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_92_pipeReg__1 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_92_pipeReg_1_0 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_92_pipeReg_1_1 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_92_REG = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_93_REG = _RAND_956[5:0];
  _RAND_957 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_93_pipeReg__0 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_93_pipeReg__1 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_93_pipeReg_1_0 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_93_pipeReg_1_1 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_93_REG = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_94_REG = _RAND_962[5:0];
  _RAND_963 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_94_pipeReg__0 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_94_pipeReg__1 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_94_pipeReg_1_0 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_94_pipeReg_1_1 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_94_REG = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_95_REG = _RAND_968[5:0];
  _RAND_969 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_95_pipeReg__0 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_95_pipeReg__1 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_95_pipeReg_1_0 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_95_pipeReg_1_1 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_95_REG = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_96_REG = _RAND_974[5:0];
  _RAND_975 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_96_pipeReg__0 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_96_pipeReg__1 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_96_pipeReg_1_0 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_96_pipeReg_1_1 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_96_REG = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_97_REG = _RAND_980[5:0];
  _RAND_981 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_97_pipeReg__0 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_97_pipeReg__1 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_97_pipeReg_1_0 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_97_pipeReg_1_1 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_97_REG = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_98_REG = _RAND_986[5:0];
  _RAND_987 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_98_pipeReg__0 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_98_pipeReg__1 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_98_pipeReg_1_0 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_98_pipeReg_1_1 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_98_REG = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_99_REG = _RAND_992[5:0];
  _RAND_993 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_99_pipeReg__0 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_99_pipeReg__1 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_99_pipeReg_1_0 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_99_pipeReg_1_1 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_99_REG = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_100_REG = _RAND_998[5:0];
  _RAND_999 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_100_pipeReg__0 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_100_pipeReg__1 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_100_pipeReg_1_0 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_100_pipeReg_1_1 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_100_REG = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_101_REG = _RAND_1004[5:0];
  _RAND_1005 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_101_pipeReg__0 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_101_pipeReg__1 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_101_pipeReg_1_0 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_101_pipeReg_1_1 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_101_REG = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_102_REG = _RAND_1010[5:0];
  _RAND_1011 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_102_pipeReg__0 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_102_pipeReg__1 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_102_pipeReg_1_0 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_102_pipeReg_1_1 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_102_REG = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_103_REG = _RAND_1016[5:0];
  _RAND_1017 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_103_pipeReg__0 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_103_pipeReg__1 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_103_pipeReg_1_0 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_103_pipeReg_1_1 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_103_REG = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_104_REG = _RAND_1022[5:0];
  _RAND_1023 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_104_pipeReg__0 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_104_pipeReg__1 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_104_pipeReg_1_0 = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_104_pipeReg_1_1 = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_104_REG = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_105_REG = _RAND_1028[5:0];
  _RAND_1029 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_105_pipeReg__0 = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_105_pipeReg__1 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_105_pipeReg_1_0 = _RAND_1031[0:0];
  _RAND_1032 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_105_pipeReg_1_1 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_105_REG = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_106_REG = _RAND_1034[5:0];
  _RAND_1035 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_106_pipeReg__0 = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_106_pipeReg__1 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_106_pipeReg_1_0 = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_106_pipeReg_1_1 = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_106_REG = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_107_REG = _RAND_1040[5:0];
  _RAND_1041 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_107_pipeReg__0 = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_107_pipeReg__1 = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_107_pipeReg_1_0 = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_107_pipeReg_1_1 = _RAND_1044[0:0];
  _RAND_1045 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_107_REG = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_108_REG = _RAND_1046[5:0];
  _RAND_1047 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_108_pipeReg__0 = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_108_pipeReg__1 = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_108_pipeReg_1_0 = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_108_pipeReg_1_1 = _RAND_1050[0:0];
  _RAND_1051 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_108_REG = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_109_REG = _RAND_1052[5:0];
  _RAND_1053 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_109_pipeReg__0 = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_109_pipeReg__1 = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_109_pipeReg_1_0 = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_109_pipeReg_1_1 = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_109_REG = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_110_REG = _RAND_1058[5:0];
  _RAND_1059 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_110_pipeReg__0 = _RAND_1059[0:0];
  _RAND_1060 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_110_pipeReg__1 = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_110_pipeReg_1_0 = _RAND_1061[0:0];
  _RAND_1062 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_110_pipeReg_1_1 = _RAND_1062[0:0];
  _RAND_1063 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_110_REG = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_111_REG = _RAND_1064[5:0];
  _RAND_1065 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_111_pipeReg__0 = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_111_pipeReg__1 = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_111_pipeReg_1_0 = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_111_pipeReg_1_1 = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_111_REG = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_112_REG = _RAND_1070[5:0];
  _RAND_1071 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_112_pipeReg__0 = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_112_pipeReg__1 = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_112_pipeReg_1_0 = _RAND_1073[0:0];
  _RAND_1074 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_112_pipeReg_1_1 = _RAND_1074[0:0];
  _RAND_1075 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_112_REG = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_113_REG = _RAND_1076[5:0];
  _RAND_1077 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_113_pipeReg__0 = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_113_pipeReg__1 = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_113_pipeReg_1_0 = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_113_pipeReg_1_1 = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_113_REG = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_114_REG = _RAND_1082[5:0];
  _RAND_1083 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_114_pipeReg__0 = _RAND_1083[0:0];
  _RAND_1084 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_114_pipeReg__1 = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_114_pipeReg_1_0 = _RAND_1085[0:0];
  _RAND_1086 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_114_pipeReg_1_1 = _RAND_1086[0:0];
  _RAND_1087 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_114_REG = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_115_REG = _RAND_1088[5:0];
  _RAND_1089 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_115_pipeReg__0 = _RAND_1089[0:0];
  _RAND_1090 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_115_pipeReg__1 = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_115_pipeReg_1_0 = _RAND_1091[0:0];
  _RAND_1092 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_115_pipeReg_1_1 = _RAND_1092[0:0];
  _RAND_1093 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_115_REG = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_116_REG = _RAND_1094[5:0];
  _RAND_1095 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_116_pipeReg__0 = _RAND_1095[0:0];
  _RAND_1096 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_116_pipeReg__1 = _RAND_1096[0:0];
  _RAND_1097 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_116_pipeReg_1_0 = _RAND_1097[0:0];
  _RAND_1098 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_116_pipeReg_1_1 = _RAND_1098[0:0];
  _RAND_1099 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_116_REG = _RAND_1099[0:0];
  _RAND_1100 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_117_REG = _RAND_1100[5:0];
  _RAND_1101 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_117_pipeReg__0 = _RAND_1101[0:0];
  _RAND_1102 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_117_pipeReg__1 = _RAND_1102[0:0];
  _RAND_1103 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_117_pipeReg_1_0 = _RAND_1103[0:0];
  _RAND_1104 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_117_pipeReg_1_1 = _RAND_1104[0:0];
  _RAND_1105 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_117_REG = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_118_REG = _RAND_1106[5:0];
  _RAND_1107 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_118_pipeReg__0 = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_118_pipeReg__1 = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_118_pipeReg_1_0 = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_118_pipeReg_1_1 = _RAND_1110[0:0];
  _RAND_1111 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_118_REG = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_119_REG = _RAND_1112[5:0];
  _RAND_1113 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_119_pipeReg__0 = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_119_pipeReg__1 = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_119_pipeReg_1_0 = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_119_pipeReg_1_1 = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_119_REG = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_120_REG = _RAND_1118[5:0];
  _RAND_1119 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_120_pipeReg__0 = _RAND_1119[0:0];
  _RAND_1120 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_120_pipeReg__1 = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_120_pipeReg_1_0 = _RAND_1121[0:0];
  _RAND_1122 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_120_pipeReg_1_1 = _RAND_1122[0:0];
  _RAND_1123 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_120_REG = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_121_REG = _RAND_1124[5:0];
  _RAND_1125 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_121_pipeReg__0 = _RAND_1125[0:0];
  _RAND_1126 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_121_pipeReg__1 = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_121_pipeReg_1_0 = _RAND_1127[0:0];
  _RAND_1128 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_121_pipeReg_1_1 = _RAND_1128[0:0];
  _RAND_1129 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_121_REG = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_122_REG = _RAND_1130[5:0];
  _RAND_1131 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_122_pipeReg__0 = _RAND_1131[0:0];
  _RAND_1132 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_122_pipeReg__1 = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_122_pipeReg_1_0 = _RAND_1133[0:0];
  _RAND_1134 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_122_pipeReg_1_1 = _RAND_1134[0:0];
  _RAND_1135 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_122_REG = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_123_REG = _RAND_1136[5:0];
  _RAND_1137 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_123_pipeReg__0 = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_123_pipeReg__1 = _RAND_1138[0:0];
  _RAND_1139 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_123_pipeReg_1_0 = _RAND_1139[0:0];
  _RAND_1140 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_123_pipeReg_1_1 = _RAND_1140[0:0];
  _RAND_1141 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_123_REG = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_124_REG = _RAND_1142[5:0];
  _RAND_1143 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_124_pipeReg__0 = _RAND_1143[0:0];
  _RAND_1144 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_124_pipeReg__1 = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_124_pipeReg_1_0 = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_124_pipeReg_1_1 = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_124_REG = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_125_REG = _RAND_1148[5:0];
  _RAND_1149 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_125_pipeReg__0 = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_125_pipeReg__1 = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_125_pipeReg_1_0 = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_125_pipeReg_1_1 = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_125_REG = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_126_REG = _RAND_1154[5:0];
  _RAND_1155 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_126_pipeReg__0 = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_126_pipeReg__1 = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_126_pipeReg_1_0 = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_126_pipeReg_1_1 = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_126_REG = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_127_REG = _RAND_1160[5:0];
  _RAND_1161 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_127_pipeReg__0 = _RAND_1161[0:0];
  _RAND_1162 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_127_pipeReg__1 = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_127_pipeReg_1_0 = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_127_pipeReg_1_1 = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_127_REG = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  pixelColorSprite = _RAND_1166[5:0];
  _RAND_1167 = {1{`RANDOM}};
  pixelColorSpriteValid = _RAND_1167[0:0];
  _RAND_1168 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_0 = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_1 = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_2 = _RAND_1170[0:0];
  _RAND_1171 = {1{`RANDOM}};
  io_vgaRed_REG = _RAND_1171[3:0];
  _RAND_1172 = {1{`RANDOM}};
  io_vgaGreen_REG = _RAND_1172[3:0];
  _RAND_1173 = {1{`RANDOM}};
  io_vgaBlue_REG = _RAND_1173[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Memory_195(
  input         clock,
  input  [7:0]  io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [27:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [7:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(8), .DATA_WIDTH(28), .LOAD_FILE("memory_init/tune_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 28'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_196(
  input         clock,
  input  [7:0]  io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [27:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [7:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(8), .DATA_WIDTH(28), .LOAD_FILE("memory_init/tune_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 28'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module SoundEngine(
  input   clock,
  input   reset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  tuneMemories_0_clock; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [7:0] tuneMemories_0_io_address; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [27:0] tuneMemories_0_io_dataRead; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire  tuneMemories_1_clock; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [7:0] tuneMemories_1_io_address; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [27:0] tuneMemories_1_io_dataRead; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  reg [11:0] durationCountReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
  reg [11:0] durationCountReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
  reg [11:0] currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
  reg [11:0] currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
  reg [7:0] nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
  reg [7:0] nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
  reg [1:0] stateReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
  reg [1:0] stateReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
  reg  newNoteLoadReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
  reg  newNoteLoadReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
  wire  durationCountRegDone_0 = durationCountReg_0 == 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 89:54]
  wire  _T_8 = tuneMemories_0_io_dataRead[27:16] != 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 111:60]
  wire [1:0] _GEN_4 = tuneMemories_0_io_dataRead[27:16] != 12'h0 ? 2'h3 : stateReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 112:23 62:25]
  wire [11:0] _GEN_6 = tuneMemories_0_io_dataRead[27:16] != 12'h0 ? tuneMemories_0_io_dataRead[27:16] :
    currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 114:30 58:32]
  wire  _T_13 = durationCountRegDone_0 & ~newNoteLoadReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:44]
  wire [7:0] _nextIndexReg_0_T_1 = nextIndexReg_0 + 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 126:46]
  wire [11:0] _GEN_10 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? tuneMemories_0_io_dataRead[27:16] :
    currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 124:30 58:32]
  wire [7:0] _GEN_12 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? _nextIndexReg_0_T_1 : nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 126:27 59:29]
  wire [7:0] _GEN_14 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? 8'h0 : _GEN_12; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 120:27]
  wire [11:0] _GEN_16 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? currDurationReg_0 : _GEN_10; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 58:32]
  wire  _GEN_17 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? 1'h0 : _T_13; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 97:23]
  wire [7:0] _GEN_22 = 2'h3 == stateReg_0 ? _GEN_14 : nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 59:29]
  wire [11:0] _GEN_24 = 2'h3 == stateReg_0 ? _GEN_16 : currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 58:32]
  wire  _GEN_25 = 2'h3 == stateReg_0 & _GEN_17; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 97:23]
  wire  durationCountRegDone_1 = durationCountReg_1 == 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 89:54]
  wire  _T_25 = tuneMemories_1_io_dataRead[27:16] != 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 111:60]
  wire [1:0] _GEN_52 = tuneMemories_1_io_dataRead[27:16] != 12'h0 ? 2'h3 : stateReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 112:23 62:25]
  wire [11:0] _GEN_54 = tuneMemories_1_io_dataRead[27:16] != 12'h0 ? tuneMemories_1_io_dataRead[27:16] :
    currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 114:30 58:32]
  wire  _T_30 = durationCountRegDone_1 & ~newNoteLoadReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:44]
  wire [7:0] _nextIndexReg_1_T_1 = nextIndexReg_1 + 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 126:46]
  wire [11:0] _GEN_58 = durationCountRegDone_1 & ~newNoteLoadReg_1 ? tuneMemories_1_io_dataRead[27:16] :
    currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 124:30 58:32]
  wire [7:0] _GEN_60 = durationCountRegDone_1 & ~newNoteLoadReg_1 ? _nextIndexReg_1_T_1 : nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 126:27 59:29]
  wire [7:0] _GEN_62 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? 8'h0 : _GEN_60; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 120:27]
  wire [11:0] _GEN_64 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? currDurationReg_1 : _GEN_58; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 58:32]
  wire  _GEN_65 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? 1'h0 : _T_30; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 97:23]
  wire [7:0] _GEN_70 = 2'h3 == stateReg_1 ? _GEN_62 : nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 59:29]
  wire [11:0] _GEN_72 = 2'h3 == stateReg_1 ? _GEN_64 : currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 58:32]
  wire  _GEN_73 = 2'h3 == stateReg_1 & _GEN_65; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 97:23]
  Memory_195 tuneMemories_0 ( // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
    .clock(tuneMemories_0_clock),
    .io_address(tuneMemories_0_io_address),
    .io_dataRead(tuneMemories_0_io_dataRead)
  );
  Memory_196 tuneMemories_1 ( // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
    .clock(tuneMemories_1_clock),
    .io_address(tuneMemories_1_io_address),
    .io_dataRead(tuneMemories_1_io_dataRead)
  );
  assign tuneMemories_0_clock = clock;
  assign tuneMemories_0_io_address = nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 72:32]
  assign tuneMemories_1_clock = clock;
  assign tuneMemories_1_io_address = nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 72:32]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
      durationCountReg_0 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
    end else if (newNoteLoadReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 84:35]
      durationCountReg_0 <= currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 85:27]
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
      durationCountReg_1 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
    end else if (newNoteLoadReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 84:35]
      durationCountReg_1 <= currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 85:27]
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
      currDurationReg_0 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
    end else if (!(2'h0 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h1 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
          currDurationReg_0 <= _GEN_6;
        end else begin
          currDurationReg_0 <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
      currDurationReg_1 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
    end else if (!(2'h0 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h1 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
          currDurationReg_1 <= _GEN_54;
        end else begin
          currDurationReg_1 <= _GEN_72;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
      nextIndexReg_0 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 102:25]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 107:25]
    end else if (!(2'h2 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= _GEN_22;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
      nextIndexReg_1 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 102:25]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 107:25]
    end else if (!(2'h2 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= _GEN_70;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
      stateReg_0 <= 2'h0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= 2'h1; // @[\\src\\main\\scala\\SoundEngine.scala 103:21]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= 2'h2; // @[\\src\\main\\scala\\SoundEngine.scala 108:21]
    end else if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= _GEN_4;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
      stateReg_1 <= 2'h0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= 2'h1; // @[\\src\\main\\scala\\SoundEngine.scala 103:21]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= 2'h2; // @[\\src\\main\\scala\\SoundEngine.scala 108:21]
    end else if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= _GEN_52;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= _T_8;
    end else begin
      newNoteLoadReg_0 <= _GEN_25;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= _T_25;
    end else begin
      newNoteLoadReg_1 <= _GEN_73;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  durationCountReg_0 = _RAND_0[11:0];
  _RAND_1 = {1{`RANDOM}};
  durationCountReg_1 = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  currDurationReg_0 = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  currDurationReg_1 = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  nextIndexReg_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  nextIndexReg_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  stateReg_0 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  stateReg_1 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  newNoteLoadReg_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  newNoteLoadReg_1 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Difficulty(
  input         clock,
  input         reset,
  input  [1:0]  io_level, // @[\\src\\main\\scala\\Difficulty.scala 5:14]
  output [26:0] io_speed, // @[\\src\\main\\scala\\Difficulty.scala 5:14]
  input         io_resetSpeed // @[\\src\\main\\scala\\Difficulty.scala 5:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [26:0] speedCnt; // @[\\src\\main\\scala\\Difficulty.scala 13:25]
  reg [26:0] frameDivider; // @[\\src\\main\\scala\\Difficulty.scala 16:29]
  wire  tick = frameDivider == 27'h196e6a; // @[\\src\\main\\scala\\Difficulty.scala 23:21]
  wire [26:0] _frameDivider_T_1 = frameDivider + 27'h1; // @[\\src\\main\\scala\\Difficulty.scala 27:34]
  wire [26:0] _speedCnt_T_1 = speedCnt + 27'h1; // @[\\src\\main\\scala\\Difficulty.scala 34:26]
  wire [21:0] timeInSeconds = speedCnt[26:5]; // @[\\src\\main\\scala\\Difficulty.scala 39:32]
  wire [18:0] scaledTime = timeInSeconds[21:3]; // @[\\src\\main\\scala\\Difficulty.scala 40:34]
  wire  _speedFactor_T = 2'h1 == io_level; // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [1:0] _speedFactor_T_1 = 2'h1 == io_level ? $signed(2'sh1) : $signed(2'sh0); // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire  _speedFactor_T_2 = 2'h2 == io_level; // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [1:0] _speedFactor_T_3 = 2'h2 == io_level ? $signed(2'sh1) : $signed(_speedFactor_T_1); // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire  _speedFactor_T_4 = 2'h3 == io_level; // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [2:0] speedFactor = 2'h3 == io_level ? $signed(3'sh2) : $signed({{1{_speedFactor_T_3[1]}},_speedFactor_T_3}); // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [20:0] _rawSpeed_T = scaledTime * 2'h3; // @[\\src\\main\\scala\\Difficulty.scala 48:37]
  wire [23:0] _rawSpeed_T_1 = $signed(_rawSpeed_T) * $signed(speedFactor); // @[\\src\\main\\scala\\Difficulty.scala 48:44]
  wire [23:0] rawSpeed = 24'sh2 + $signed(_rawSpeed_T_1); // @[\\src\\main\\scala\\Difficulty.scala 48:22]
  wire [4:0] _speedCap_T_1 = _speedFactor_T ? $signed(5'shc) : $signed(5'sha); // @[\\src\\main\\scala\\Difficulty.scala 50:43]
  wire [5:0] _speedCap_T_3 = _speedFactor_T_2 ? $signed(6'sh10) : $signed({{1{_speedCap_T_1[4]}},_speedCap_T_1}); // @[\\src\\main\\scala\\Difficulty.scala 50:43]
  wire [5:0] speedCap = _speedFactor_T_4 ? $signed(6'sh16) : $signed(_speedCap_T_3); // @[\\src\\main\\scala\\Difficulty.scala 50:43]
  wire [23:0] _GEN_4 = {{18{speedCap[5]}},speedCap}; // @[\\src\\main\\scala\\Difficulty.scala 55:28]
  wire [23:0] _io_speed_T_1 = $signed(rawSpeed) > $signed(_GEN_4) ? $signed({{18{speedCap[5]}},speedCap}) : $signed(
    rawSpeed); // @[\\src\\main\\scala\\Difficulty.scala 55:18]
  assign io_speed = {{3{_io_speed_T_1[23]}},_io_speed_T_1}; // @[\\src\\main\\scala\\Difficulty.scala 55:12]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\Difficulty.scala 13:25]
      speedCnt <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 13:25]
    end else if (io_resetSpeed) begin // @[\\src\\main\\scala\\Difficulty.scala 31:23]
      speedCnt <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 32:14]
    end else if (tick) begin // @[\\src\\main\\scala\\Difficulty.scala 33:20]
      speedCnt <= _speedCnt_T_1; // @[\\src\\main\\scala\\Difficulty.scala 34:14]
    end
    if (reset) begin // @[\\src\\main\\scala\\Difficulty.scala 16:29]
      frameDivider <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 16:29]
    end else if (tick) begin // @[\\src\\main\\scala\\Difficulty.scala 23:37]
      frameDivider <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 24:18]
    end else begin
      frameDivider <= _frameDivider_T_1; // @[\\src\\main\\scala\\Difficulty.scala 27:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  speedCnt = _RAND_0[26:0];
  _RAND_1 = {1{`RANDOM}};
  frameDivider = _RAND_1[26:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LFSR(
  input        clock,
  input        reset,
  output [9:0] io_out_0, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_1, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_2, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_3, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_4, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_5, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_6, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_7, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_8, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_9, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_10, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_11, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_12, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_13, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_14, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_15, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_16, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_17, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_18, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_19, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_20, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_21, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_22, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_23, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_24, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_25, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_26, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_27, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_28, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_29 // @[\\src\\main\\scala\\LFSR.scala 5:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] reg_; // @[\\src\\main\\scala\\LFSR.scala 10:20]
  wire  feedback = reg_[63] ^ reg_[62] ^ reg_[60] ^ reg_[59]; // @[\\src\\main\\scala\\LFSR.scala 13:46]
  wire [63:0] _reg_T_1 = {reg_[62:0],feedback}; // @[\\src\\main\\scala\\LFSR.scala 16:13]
  wire [8:0] current_output = reg_[17:9]; // @[\\src\\main\\scala\\LFSR.scala 19:27]
  reg [9:0] history_0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_1; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_2; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_3; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_4; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_5; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_6; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_7; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_8; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_9; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_10; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_11; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_12; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_13; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_14; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_15; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_16; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_17; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_18; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_19; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_20; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_21; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_22; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_23; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_24; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_25; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_26; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_27; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_28; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_29; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  assign io_out_0 = history_0; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_1 = history_1; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_2 = history_2; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_3 = history_3; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_4 = history_4; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_5 = history_5; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_6 = history_6; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_7 = history_7; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_8 = history_8; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_9 = history_9; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_10 = history_10; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_11 = history_11; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_12 = history_12; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_13 = history_13; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_14 = history_14; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_15 = history_15; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_16 = history_16; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_17 = history_17; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_18 = history_18; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_19 = history_19; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_20 = history_20; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_21 = history_21; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_22 = history_22; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_23 = history_23; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_24 = history_24; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_25 = history_25; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_26 = history_26; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_27 = history_27; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_28 = history_28; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_29 = history_29; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 10:20]
      reg_ <= 64'h123456789abcdef; // @[\\src\\main\\scala\\LFSR.scala 10:20]
    end else begin
      reg_ <= _reg_T_1; // @[\\src\\main\\scala\\LFSR.scala 16:7]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_0 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_0 <= history_1; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_1 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_1 <= history_2; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_2 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_2 <= history_3; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_3 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_3 <= history_4; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_4 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_4 <= history_5; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_5 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_5 <= history_6; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_6 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_6 <= history_7; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_7 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_7 <= history_8; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_8 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_8 <= history_9; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_9 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_9 <= history_10; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_10 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_10 <= history_11; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_11 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_11 <= history_12; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_12 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_12 <= history_13; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_13 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_13 <= history_14; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_14 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_14 <= history_15; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_15 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_15 <= history_16; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_16 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_16 <= history_17; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_17 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_17 <= history_18; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_18 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_18 <= history_19; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_19 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_19 <= history_20; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_20 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_20 <= history_21; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_21 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_21 <= history_22; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_22 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_22 <= history_23; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_23 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_23 <= history_24; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_24 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_24 <= history_25; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_25 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_25 <= history_26; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_26 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_26 <= history_27; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_27 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_27 <= history_28; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_28 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_28 <= history_29; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_29 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_29 <= {{1'd0}, current_output}; // @[\\src\\main\\scala\\LFSR.scala 28:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_ = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  history_0 = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  history_1 = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  history_2 = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  history_3 = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  history_4 = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  history_5 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  history_6 = _RAND_7[9:0];
  _RAND_8 = {1{`RANDOM}};
  history_7 = _RAND_8[9:0];
  _RAND_9 = {1{`RANDOM}};
  history_8 = _RAND_9[9:0];
  _RAND_10 = {1{`RANDOM}};
  history_9 = _RAND_10[9:0];
  _RAND_11 = {1{`RANDOM}};
  history_10 = _RAND_11[9:0];
  _RAND_12 = {1{`RANDOM}};
  history_11 = _RAND_12[9:0];
  _RAND_13 = {1{`RANDOM}};
  history_12 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  history_13 = _RAND_14[9:0];
  _RAND_15 = {1{`RANDOM}};
  history_14 = _RAND_15[9:0];
  _RAND_16 = {1{`RANDOM}};
  history_15 = _RAND_16[9:0];
  _RAND_17 = {1{`RANDOM}};
  history_16 = _RAND_17[9:0];
  _RAND_18 = {1{`RANDOM}};
  history_17 = _RAND_18[9:0];
  _RAND_19 = {1{`RANDOM}};
  history_18 = _RAND_19[9:0];
  _RAND_20 = {1{`RANDOM}};
  history_19 = _RAND_20[9:0];
  _RAND_21 = {1{`RANDOM}};
  history_20 = _RAND_21[9:0];
  _RAND_22 = {1{`RANDOM}};
  history_21 = _RAND_22[9:0];
  _RAND_23 = {1{`RANDOM}};
  history_22 = _RAND_23[9:0];
  _RAND_24 = {1{`RANDOM}};
  history_23 = _RAND_24[9:0];
  _RAND_25 = {1{`RANDOM}};
  history_24 = _RAND_25[9:0];
  _RAND_26 = {1{`RANDOM}};
  history_25 = _RAND_26[9:0];
  _RAND_27 = {1{`RANDOM}};
  history_26 = _RAND_27[9:0];
  _RAND_28 = {1{`RANDOM}};
  history_27 = _RAND_28[9:0];
  _RAND_29 = {1{`RANDOM}};
  history_28 = _RAND_29[9:0];
  _RAND_30 = {1{`RANDOM}};
  history_29 = _RAND_30[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GameLogic(
  input         clock,
  input         reset,
  input         io_btnC, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnU, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnL, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnR, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnD, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_3, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_7, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_8, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_9, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_10, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_11, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_12, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_13, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_14, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_46, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_47, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_48, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_49, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_50, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_51, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_52, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_53, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_54, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_55, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_56, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_57, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_61, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_62, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_63, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_3, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_7, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_8, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_9, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_10, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_11, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_12, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_13, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_14, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_46, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_47, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_48, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_49, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_50, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_51, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_52, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_53, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_54, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_55, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_56, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_57, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_61, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_62, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_63, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_3, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_4, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_5, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_6, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_7, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_8, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_9, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_10, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_11, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_12, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_13, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_14, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_15, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_46, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_47, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_48, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_49, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_50, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_51, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_52, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_53, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_54, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_55, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_56, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_57, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_61, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_62, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_63, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_64, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_65, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_66, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_67, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_68, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_69, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_70, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_71, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_72, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_73, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_74, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_75, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_76, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_77, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_78, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_79, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_80, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_81, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_82, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_83, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_84, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_85, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_86, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_87, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_88, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_89, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_90, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_91, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_92, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_93, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_94, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_95, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_96, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_97, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_98, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_99, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_viewBoxX, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [8:0]  io_viewBoxY, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_newFrame, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_frameUpdateDone // @[\\src\\main\\scala\\GameLogic.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
`endif // RANDOMIZE_REG_INIT
  wire  difficulty_clock; // @[\\src\\main\\scala\\GameLogic.scala 217:26]
  wire  difficulty_reset; // @[\\src\\main\\scala\\GameLogic.scala 217:26]
  wire [1:0] difficulty_io_level; // @[\\src\\main\\scala\\GameLogic.scala 217:26]
  wire [26:0] difficulty_io_speed; // @[\\src\\main\\scala\\GameLogic.scala 217:26]
  wire  difficulty_io_resetSpeed; // @[\\src\\main\\scala\\GameLogic.scala 217:26]
  wire  lfsr_clock; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire  lfsr_reset; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_0; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_1; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_2; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_3; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_4; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_5; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_6; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_7; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_8; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_9; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_10; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_11; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_12; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_13; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_14; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_15; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_16; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_17; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_18; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_19; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_20; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_21; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_22; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_23; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_24; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_25; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_26; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_27; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_28; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  wire [9:0] lfsr_io_out_29; // @[\\src\\main\\scala\\GameLogic.scala 259:20]
  reg [2:0] stateReg; // @[\\src\\main\\scala\\GameLogic.scala 113:25]
  reg [10:0] spriteXRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [9:0] spriteYRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg  spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_64; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_65; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_66; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_67; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_68; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_69; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_70; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_71; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_72; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_73; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_74; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_75; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_76; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_77; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_78; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_79; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_80; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_81; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_82; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_83; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_84; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_85; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_86; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_87; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_88; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_89; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_90; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_91; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_92; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_93; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_94; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_95; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_96; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_97; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_98; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_99; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  initializePositions; // @[\\src\\main\\scala\\GameLogic.scala 130:36]
  wire [10:0] _GEN_0 = initializePositions ? $signed(11'sh140) : $signed(spriteXRegs_3); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_1 = initializePositions ? $signed(10'shf0) : $signed(spriteYRegs_3); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_14 = initializePositions ? $signed(11'sh140) : $signed(spriteXRegs_13); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_15 = initializePositions ? $signed(10'shf0) : $signed(spriteYRegs_13); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_16 = initializePositions ? $signed(11'sh260) : $signed(spriteXRegs_14); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_17 = initializePositions ? $signed(10'shf0) : $signed(spriteYRegs_14); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_18 = initializePositions ? $signed(11'sh168) : $signed(spriteXRegs_16); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_19 = initializePositions ? $signed(10'sh14) : $signed(spriteYRegs_16); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_20 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_17); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_21 = initializePositions ? $signed(10'sh32) : $signed(spriteYRegs_17); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_22 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_18); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_23 = initializePositions ? $signed(10'sh50) : $signed(spriteYRegs_18); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_24 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_19); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_25 = initializePositions ? $signed(10'sh6e) : $signed(spriteYRegs_19); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_26 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_20); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_27 = initializePositions ? $signed(10'sh8c) : $signed(spriteYRegs_20); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_28 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_21); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_29 = initializePositions ? $signed(10'shaa) : $signed(spriteYRegs_21); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_30 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_22); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_31 = initializePositions ? $signed(10'shc8) : $signed(spriteYRegs_22); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_32 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_23); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_33 = initializePositions ? $signed(10'she6) : $signed(spriteYRegs_23); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_34 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_24); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_35 = initializePositions ? $signed(10'sh104) : $signed(spriteYRegs_24); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_36 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_25); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_37 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_25); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_38 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_26); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_39 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_26); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_40 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_27); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_41 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_27); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_42 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_28); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_43 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_28); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_44 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_29); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_45 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_29); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_46 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_30); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_47 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_30); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_48 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_31); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_49 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_31); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_50 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_32); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_51 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_32); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_52 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_33); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_53 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_33); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_54 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_34); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_55 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_34); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_56 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_35); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_57 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_35); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_58 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_36); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_59 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_36); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_60 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_37); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_61 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_37); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_62 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_38); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_63 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_38); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_64 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_39); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_65 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_39); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_66 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_40); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_67 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_40); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_68 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_41); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_69 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_41); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_70 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_42); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_71 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_42); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_72 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_43); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_73 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_43); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_74 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_44); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_75 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_44); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_76 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_45); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_77 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_45); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_102 = initializePositions ? $signed(11'sh140) : $signed(spriteXRegs_58); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_103 = initializePositions ? $signed(10'sh14) : $signed(spriteYRegs_58); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_104 = initializePositions ? $signed(11'sh1f4) : $signed(spriteXRegs_59); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_105 = initializePositions ? $signed(10'sh46) : $signed(spriteYRegs_59); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire [10:0] _GEN_106 = initializePositions ? $signed(11'sh96) : $signed(spriteXRegs_60); // @[\\src\\main\\scala\\GameLogic.scala 131:29 169:23 121:28]
  wire [9:0] _GEN_107 = initializePositions ? $signed(10'sh64) : $signed(spriteYRegs_60); // @[\\src\\main\\scala\\GameLogic.scala 131:29 170:23 122:28]
  wire  _GEN_186 = initializePositions ? 1'h0 : initializePositions; // @[\\src\\main\\scala\\GameLogic.scala 131:29 172:25 130:36]
  reg  sprite58ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 176:42]
  reg  sprite58ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 177:40]
  reg  sprite59ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 178:42]
  reg  sprite59ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 179:40]
  reg  sprite60ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 180:42]
  reg  sprite60ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 181:40]
  reg [9:0] viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 209:28]
  reg [8:0] viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 210:28]
  reg [1:0] lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 219:23]
  reg [2:0] livesReg; // @[\\src\\main\\scala\\GameLogic.scala 231:25]
  reg [9:0] extraLifeCnt; // @[\\src\\main\\scala\\GameLogic.scala 234:29]
  reg  gameOverReturnPressed; // @[\\src\\main\\scala\\GameLogic.scala 237:38]
  reg [7:0] spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 243:34]
  reg [5:0] nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 244:34]
  reg [9:0] starCnt; // @[\\src\\main\\scala\\GameLogic.scala 247:24]
  reg  collisionDetected; // @[\\src\\main\\scala\\GameLogic.scala 250:34]
  reg [7:0] blinkCounter; // @[\\src\\main\\scala\\GameLogic.scala 251:29]
  reg [1:0] blinkTimes; // @[\\src\\main\\scala\\GameLogic.scala 252:27]
  reg  isBlinking; // @[\\src\\main\\scala\\GameLogic.scala 253:27]
  wire  _T = lvlReg != 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 262:15]
  wire  _T_1 = livesReg == 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 263:19]
  wire  _T_2 = livesReg == 3'h2; // @[\\src\\main\\scala\\GameLogic.scala 267:25]
  wire  _T_3 = livesReg == 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 271:25]
  wire  _GEN_189 = livesReg == 3'h2 | _T_3; // @[\\src\\main\\scala\\GameLogic.scala 267:34 268:29]
  wire  _GEN_192 = livesReg == 3'h3 | _GEN_189; // @[\\src\\main\\scala\\GameLogic.scala 263:28 264:29]
  wire  _GEN_193 = livesReg == 3'h3 | _T_2; // @[\\src\\main\\scala\\GameLogic.scala 263:28 265:29]
  wire  _GEN_195 = lvlReg != 2'h0 & _GEN_192; // @[\\src\\main\\scala\\GameLogic.scala 262:24 281:27]
  wire  _GEN_196 = lvlReg != 2'h0 & _GEN_193; // @[\\src\\main\\scala\\GameLogic.scala 262:24 282:27]
  wire  _GEN_197 = lvlReg != 2'h0 & _T_1; // @[\\src\\main\\scala\\GameLogic.scala 262:24 283:27]
  wire  _T_5 = livesReg == 3'h0; // @[\\src\\main\\scala\\GameLogic.scala 353:29]
  wire [2:0] _GEN_198 = livesReg == 3'h0 ? 3'h6 : 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 353:38 354:20 356:20]
  wire  _GEN_210 = gameOverReturnPressed | _GEN_186; // @[\\src\\main\\scala\\GameLogic.scala 302:25 349:37]
  wire  _GEN_211 = gameOverReturnPressed | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 305:26 125:34 349:37]
  wire  _GEN_268 = io_newFrame ? _GEN_210 : _GEN_186; // @[\\src\\main\\scala\\GameLogic.scala 348:25]
  wire [9:0] _spriteYRegs_16_T_2 = 10'h64 + lfsr_io_out_0; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_201 = {{16{spriteXRegs_16[10]}},spriteXRegs_16}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_16_T_2 = $signed(_GEN_201) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_315 = spriteVisibleRegs_16 ? $signed(_spriteXRegs_16_T_2) : $signed({{16{_GEN_18[10]}},_GEN_18}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_316 = $signed(spriteXRegs_16) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_315); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_317 = $signed(spriteXRegs_16) >= 11'sh280 ? $signed(_spriteYRegs_16_T_2) : $signed(_GEN_19); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_318 = $signed(spriteXRegs_16) >= 11'sh280 ? lfsr_io_out_10[0] : spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_319 = ~spriteScaleTypeRegs_0 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [9:0] _spriteYRegs_17_T_2 = 10'h64 + lfsr_io_out_1; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_259 = {{16{spriteXRegs_17[10]}},spriteXRegs_17}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_17_T_2 = $signed(_GEN_259) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_320 = spriteVisibleRegs_17 ? $signed(_spriteXRegs_17_T_2) : $signed({{16{_GEN_20[10]}},_GEN_20}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_321 = $signed(spriteXRegs_17) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_320); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_322 = $signed(spriteXRegs_17) >= 11'sh280 ? $signed(_spriteYRegs_17_T_2) : $signed(_GEN_21); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_323 = $signed(spriteXRegs_17) >= 11'sh280 ? lfsr_io_out_11[0] : spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_324 = ~spriteScaleTypeRegs_1 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [9:0] _spriteYRegs_18_T_2 = 10'h64 + lfsr_io_out_2; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_605 = {{16{spriteXRegs_18[10]}},spriteXRegs_18}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_18_T_2 = $signed(_GEN_605) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_325 = spriteVisibleRegs_18 ? $signed(_spriteXRegs_18_T_2) : $signed({{16{_GEN_22[10]}},_GEN_22}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_326 = $signed(spriteXRegs_18) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_325); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_327 = $signed(spriteXRegs_18) >= 11'sh280 ? $signed(_spriteYRegs_18_T_2) : $signed(_GEN_23); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_328 = $signed(spriteXRegs_18) >= 11'sh280 ? lfsr_io_out_12[0] : spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_329 = ~spriteScaleTypeRegs_2 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [9:0] _spriteYRegs_19_T_2 = 10'h64 + lfsr_io_out_3; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_606 = {{16{spriteXRegs_19[10]}},spriteXRegs_19}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_19_T_2 = $signed(_GEN_606) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_330 = spriteVisibleRegs_19 ? $signed(_spriteXRegs_19_T_2) : $signed({{16{_GEN_24[10]}},_GEN_24}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_331 = $signed(spriteXRegs_19) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_330); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_332 = $signed(spriteXRegs_19) >= 11'sh280 ? $signed(_spriteYRegs_19_T_2) : $signed(_GEN_25); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_333 = $signed(spriteXRegs_19) >= 11'sh280 ? lfsr_io_out_13[0] : spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_334 = ~spriteScaleTypeRegs_3 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [9:0] _spriteYRegs_20_T_2 = 10'h64 + lfsr_io_out_4; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_607 = {{16{spriteXRegs_20[10]}},spriteXRegs_20}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_20_T_2 = $signed(_GEN_607) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_335 = spriteVisibleRegs_20 ? $signed(_spriteXRegs_20_T_2) : $signed({{16{_GEN_26[10]}},_GEN_26}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_336 = $signed(spriteXRegs_20) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_335); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_337 = $signed(spriteXRegs_20) >= 11'sh280 ? $signed(_spriteYRegs_20_T_2) : $signed(_GEN_27); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_338 = $signed(spriteXRegs_20) >= 11'sh280 ? lfsr_io_out_14[0] : spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_339 = ~spriteScaleTypeRegs_4 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [9:0] _spriteYRegs_21_T_2 = 10'h64 + lfsr_io_out_5; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_663 = {{16{spriteXRegs_21[10]}},spriteXRegs_21}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_21_T_2 = $signed(_GEN_663) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_340 = spriteVisibleRegs_21 ? $signed(_spriteXRegs_21_T_2) : $signed({{16{_GEN_28[10]}},_GEN_28}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_341 = $signed(spriteXRegs_21) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_340); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_342 = $signed(spriteXRegs_21) >= 11'sh280 ? $signed(_spriteYRegs_21_T_2) : $signed(_GEN_29); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_343 = $signed(spriteXRegs_21) >= 11'sh280 ? lfsr_io_out_15[0] : spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_344 = ~spriteScaleTypeRegs_5 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [9:0] _spriteYRegs_22_T_2 = 10'h64 + lfsr_io_out_6; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_664 = {{16{spriteXRegs_22[10]}},spriteXRegs_22}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_22_T_2 = $signed(_GEN_664) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_345 = spriteVisibleRegs_22 ? $signed(_spriteXRegs_22_T_2) : $signed({{16{_GEN_30[10]}},_GEN_30}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_346 = $signed(spriteXRegs_22) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_345); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_347 = $signed(spriteXRegs_22) >= 11'sh280 ? $signed(_spriteYRegs_22_T_2) : $signed(_GEN_31); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_348 = $signed(spriteXRegs_22) >= 11'sh280 ? lfsr_io_out_16[0] : spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_349 = ~spriteScaleTypeRegs_6 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [9:0] _spriteYRegs_23_T_2 = 10'h64 + lfsr_io_out_7; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_665 = {{16{spriteXRegs_23[10]}},spriteXRegs_23}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_23_T_2 = $signed(_GEN_665) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_350 = spriteVisibleRegs_23 ? $signed(_spriteXRegs_23_T_2) : $signed({{16{_GEN_32[10]}},_GEN_32}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_351 = $signed(spriteXRegs_23) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_350); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_352 = $signed(spriteXRegs_23) >= 11'sh280 ? $signed(_spriteYRegs_23_T_2) : $signed(_GEN_33); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_353 = $signed(spriteXRegs_23) >= 11'sh280 ? lfsr_io_out_17[0] : spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_354 = ~spriteScaleTypeRegs_7 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [9:0] _spriteYRegs_24_T_2 = 10'h64 + lfsr_io_out_8; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_706 = {{16{spriteXRegs_24[10]}},spriteXRegs_24}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_24_T_2 = $signed(_GEN_706) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_355 = spriteVisibleRegs_24 ? $signed(_spriteXRegs_24_T_2) : $signed({{16{_GEN_34[10]}},_GEN_34}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_356 = $signed(spriteXRegs_24) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_355); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_357 = $signed(spriteXRegs_24) >= 11'sh280 ? $signed(_spriteYRegs_24_T_2) : $signed(_GEN_35); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_358 = $signed(spriteXRegs_24) >= 11'sh280 ? lfsr_io_out_18[0] : spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_359 = ~spriteScaleTypeRegs_8 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [9:0] _spriteYRegs_25_T_2 = 10'h64 + lfsr_io_out_9; // @[\\src\\main\\scala\\GameLogic.scala 377:63]
  wire [26:0] _GEN_707 = {{16{spriteXRegs_25[10]}},spriteXRegs_25}; // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _spriteXRegs_25_T_2 = $signed(_GEN_707) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 382:46]
  wire [26:0] _GEN_360 = spriteVisibleRegs_25 ? $signed(_spriteXRegs_25_T_2) : $signed({{16{_GEN_36[10]}},_GEN_36}); // @[\\src\\main\\scala\\GameLogic.scala 381:44 382:28]
  wire [26:0] _GEN_361 = $signed(spriteXRegs_25) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_360); // @[\\src\\main\\scala\\GameLogic.scala 375:41 376:28]
  wire [9:0] _GEN_362 = $signed(spriteXRegs_25) >= 11'sh280 ? $signed(_spriteYRegs_25_T_2) : $signed(_GEN_37); // @[\\src\\main\\scala\\GameLogic.scala 375:41 377:28]
  wire  _GEN_363 = $signed(spriteXRegs_25) >= 11'sh280 ? lfsr_io_out_19[0] : spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 126:36 375:41 379:40]
  wire  _GEN_364 = ~spriteScaleTypeRegs_9 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 386:52 387:43 390:43]
  wire [26:0] _GEN_708 = {{16{spriteXRegs_26[10]}},spriteXRegs_26}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_26_T_2 = $signed(_GEN_708) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_365 = spriteVisibleRegs_26 ? $signed(_spriteXRegs_26_T_2) : $signed({{16{_GEN_38[10]}},_GEN_38}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_366 = $signed(spriteXRegs_26) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_365); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_367 = $signed(spriteXRegs_26) >= 11'sh280 ? $signed(_spriteYRegs_16_T_2) : $signed(_GEN_39); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_368 = $signed(spriteXRegs_26) >= 11'sh280 ? lfsr_io_out_10[0] : _GEN_318; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [26:0] _GEN_764 = {{16{spriteXRegs_27[10]}},spriteXRegs_27}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_27_T_2 = $signed(_GEN_764) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_370 = spriteVisibleRegs_27 ? $signed(_spriteXRegs_27_T_2) : $signed({{16{_GEN_40[10]}},_GEN_40}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_371 = $signed(spriteXRegs_27) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_370); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_372 = $signed(spriteXRegs_27) >= 11'sh280 ? $signed(_spriteYRegs_17_T_2) : $signed(_GEN_41); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_373 = $signed(spriteXRegs_27) >= 11'sh280 ? lfsr_io_out_11[0] : _GEN_323; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [26:0] _GEN_765 = {{16{spriteXRegs_28[10]}},spriteXRegs_28}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_28_T_2 = $signed(_GEN_765) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_375 = spriteVisibleRegs_28 ? $signed(_spriteXRegs_28_T_2) : $signed({{16{_GEN_42[10]}},_GEN_42}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_376 = $signed(spriteXRegs_28) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_375); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_377 = $signed(spriteXRegs_28) >= 11'sh280 ? $signed(_spriteYRegs_18_T_2) : $signed(_GEN_43); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_378 = $signed(spriteXRegs_28) >= 11'sh280 ? lfsr_io_out_12[0] : _GEN_328; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [26:0] _GEN_766 = {{16{spriteXRegs_29[10]}},spriteXRegs_29}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_29_T_2 = $signed(_GEN_766) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_380 = spriteVisibleRegs_29 ? $signed(_spriteXRegs_29_T_2) : $signed({{16{_GEN_44[10]}},_GEN_44}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_381 = $signed(spriteXRegs_29) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_380); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_382 = $signed(spriteXRegs_29) >= 11'sh280 ? $signed(_spriteYRegs_19_T_2) : $signed(_GEN_45); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_383 = $signed(spriteXRegs_29) >= 11'sh280 ? lfsr_io_out_13[0] : _GEN_333; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [26:0] _GEN_808 = {{16{spriteXRegs_30[10]}},spriteXRegs_30}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_30_T_2 = $signed(_GEN_808) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_385 = spriteVisibleRegs_30 ? $signed(_spriteXRegs_30_T_2) : $signed({{16{_GEN_46[10]}},_GEN_46}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_386 = $signed(spriteXRegs_30) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_385); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_387 = $signed(spriteXRegs_30) >= 11'sh280 ? $signed(_spriteYRegs_20_T_2) : $signed(_GEN_47); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_388 = $signed(spriteXRegs_30) >= 11'sh280 ? lfsr_io_out_14[0] : _GEN_338; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [26:0] _GEN_809 = {{16{spriteXRegs_31[10]}},spriteXRegs_31}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_31_T_2 = $signed(_GEN_809) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_390 = spriteVisibleRegs_31 ? $signed(_spriteXRegs_31_T_2) : $signed({{16{_GEN_48[10]}},_GEN_48}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_391 = $signed(spriteXRegs_31) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_390); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_392 = $signed(spriteXRegs_31) >= 11'sh280 ? $signed(_spriteYRegs_21_T_2) : $signed(_GEN_49); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_393 = $signed(spriteXRegs_31) >= 11'sh280 ? lfsr_io_out_15[0] : _GEN_343; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [26:0] _GEN_810 = {{16{spriteXRegs_32[10]}},spriteXRegs_32}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_32_T_2 = $signed(_GEN_810) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_395 = spriteVisibleRegs_32 ? $signed(_spriteXRegs_32_T_2) : $signed({{16{_GEN_50[10]}},_GEN_50}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_396 = $signed(spriteXRegs_32) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_395); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_397 = $signed(spriteXRegs_32) >= 11'sh280 ? $signed(_spriteYRegs_22_T_2) : $signed(_GEN_51); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_398 = $signed(spriteXRegs_32) >= 11'sh280 ? lfsr_io_out_16[0] : _GEN_348; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [26:0] _GEN_866 = {{16{spriteXRegs_33[10]}},spriteXRegs_33}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_33_T_2 = $signed(_GEN_866) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_400 = spriteVisibleRegs_33 ? $signed(_spriteXRegs_33_T_2) : $signed({{16{_GEN_52[10]}},_GEN_52}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_401 = $signed(spriteXRegs_33) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_400); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_402 = $signed(spriteXRegs_33) >= 11'sh280 ? $signed(_spriteYRegs_23_T_2) : $signed(_GEN_53); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_403 = $signed(spriteXRegs_33) >= 11'sh280 ? lfsr_io_out_17[0] : _GEN_353; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [26:0] _GEN_867 = {{16{spriteXRegs_34[10]}},spriteXRegs_34}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_34_T_2 = $signed(_GEN_867) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_405 = spriteVisibleRegs_34 ? $signed(_spriteXRegs_34_T_2) : $signed({{16{_GEN_54[10]}},_GEN_54}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_406 = $signed(spriteXRegs_34) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_405); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_407 = $signed(spriteXRegs_34) >= 11'sh280 ? $signed(_spriteYRegs_24_T_2) : $signed(_GEN_55); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_408 = $signed(spriteXRegs_34) >= 11'sh280 ? lfsr_io_out_18[0] : _GEN_358; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [26:0] _GEN_868 = {{16{spriteXRegs_35[10]}},spriteXRegs_35}; // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _spriteXRegs_35_T_2 = $signed(_GEN_868) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 405:46]
  wire [26:0] _GEN_410 = spriteVisibleRegs_35 ? $signed(_spriteXRegs_35_T_2) : $signed({{16{_GEN_56[10]}},_GEN_56}); // @[\\src\\main\\scala\\GameLogic.scala 404:44 405:28]
  wire [26:0] _GEN_411 = $signed(spriteXRegs_35) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_410); // @[\\src\\main\\scala\\GameLogic.scala 398:41 399:28]
  wire [9:0] _GEN_412 = $signed(spriteXRegs_35) >= 11'sh280 ? $signed(_spriteYRegs_25_T_2) : $signed(_GEN_57); // @[\\src\\main\\scala\\GameLogic.scala 398:41 400:28]
  wire  _GEN_413 = $signed(spriteXRegs_35) >= 11'sh280 ? lfsr_io_out_19[0] : _GEN_363; // @[\\src\\main\\scala\\GameLogic.scala 398:41 402:40]
  wire [9:0] _spriteYRegs_36_T_2 = 10'h64 + lfsr_io_out_20; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_909 = {{16{spriteXRegs_36[10]}},spriteXRegs_36}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_36_T_2 = $signed(_GEN_909) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_415 = spriteVisibleRegs_36 ? $signed(_spriteXRegs_36_T_2) : $signed({{16{_GEN_58[10]}},_GEN_58}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_416 = $signed(spriteXRegs_36) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_415); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_417 = $signed(spriteXRegs_36) >= 11'sh280 ? $signed(_spriteYRegs_36_T_2) : $signed(_GEN_59); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_418 = $signed(spriteXRegs_36) >= 11'sh280 ? lfsr_io_out_10[0] : _GEN_368; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _spriteYRegs_37_T_2 = 10'h64 + lfsr_io_out_21; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_910 = {{16{spriteXRegs_37[10]}},spriteXRegs_37}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_37_T_2 = $signed(_GEN_910) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_420 = spriteVisibleRegs_37 ? $signed(_spriteXRegs_37_T_2) : $signed({{16{_GEN_60[10]}},_GEN_60}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_421 = $signed(spriteXRegs_37) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_420); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_422 = $signed(spriteXRegs_37) >= 11'sh280 ? $signed(_spriteYRegs_37_T_2) : $signed(_GEN_61); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_423 = $signed(spriteXRegs_37) >= 11'sh280 ? lfsr_io_out_11[0] : _GEN_373; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _spriteYRegs_38_T_2 = 10'h64 + lfsr_io_out_22; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_911 = {{16{spriteXRegs_38[10]}},spriteXRegs_38}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_38_T_2 = $signed(_GEN_911) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_425 = spriteVisibleRegs_38 ? $signed(_spriteXRegs_38_T_2) : $signed({{16{_GEN_62[10]}},_GEN_62}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_426 = $signed(spriteXRegs_38) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_425); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_427 = $signed(spriteXRegs_38) >= 11'sh280 ? $signed(_spriteYRegs_38_T_2) : $signed(_GEN_63); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_428 = $signed(spriteXRegs_38) >= 11'sh280 ? lfsr_io_out_12[0] : _GEN_378; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _spriteYRegs_39_T_2 = 10'h64 + lfsr_io_out_23; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_967 = {{16{spriteXRegs_39[10]}},spriteXRegs_39}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_39_T_2 = $signed(_GEN_967) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_430 = spriteVisibleRegs_39 ? $signed(_spriteXRegs_39_T_2) : $signed({{16{_GEN_64[10]}},_GEN_64}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_431 = $signed(spriteXRegs_39) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_430); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_432 = $signed(spriteXRegs_39) >= 11'sh280 ? $signed(_spriteYRegs_39_T_2) : $signed(_GEN_65); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_433 = $signed(spriteXRegs_39) >= 11'sh280 ? lfsr_io_out_13[0] : _GEN_383; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _spriteYRegs_40_T_2 = 10'h64 + lfsr_io_out_24; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_968 = {{16{spriteXRegs_40[10]}},spriteXRegs_40}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_40_T_2 = $signed(_GEN_968) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_435 = spriteVisibleRegs_40 ? $signed(_spriteXRegs_40_T_2) : $signed({{16{_GEN_66[10]}},_GEN_66}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_436 = $signed(spriteXRegs_40) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_435); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_437 = $signed(spriteXRegs_40) >= 11'sh280 ? $signed(_spriteYRegs_40_T_2) : $signed(_GEN_67); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_438 = $signed(spriteXRegs_40) >= 11'sh280 ? lfsr_io_out_14[0] : _GEN_388; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _spriteYRegs_41_T_2 = 10'h64 + lfsr_io_out_25; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_969 = {{16{spriteXRegs_41[10]}},spriteXRegs_41}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_41_T_2 = $signed(_GEN_969) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_440 = spriteVisibleRegs_41 ? $signed(_spriteXRegs_41_T_2) : $signed({{16{_GEN_68[10]}},_GEN_68}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_441 = $signed(spriteXRegs_41) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_440); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_442 = $signed(spriteXRegs_41) >= 11'sh280 ? $signed(_spriteYRegs_41_T_2) : $signed(_GEN_69); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_443 = $signed(spriteXRegs_41) >= 11'sh280 ? lfsr_io_out_15[0] : _GEN_393; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _spriteYRegs_42_T_2 = 10'h64 + lfsr_io_out_26; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_1011 = {{16{spriteXRegs_42[10]}},spriteXRegs_42}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_42_T_2 = $signed(_GEN_1011) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_445 = spriteVisibleRegs_42 ? $signed(_spriteXRegs_42_T_2) : $signed({{16{_GEN_70[10]}},_GEN_70}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_446 = $signed(spriteXRegs_42) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_445); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_447 = $signed(spriteXRegs_42) >= 11'sh280 ? $signed(_spriteYRegs_42_T_2) : $signed(_GEN_71); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_448 = $signed(spriteXRegs_42) >= 11'sh280 ? lfsr_io_out_16[0] : _GEN_398; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _spriteYRegs_43_T_2 = 10'h64 + lfsr_io_out_27; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_1012 = {{16{spriteXRegs_43[10]}},spriteXRegs_43}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_43_T_2 = $signed(_GEN_1012) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_450 = spriteVisibleRegs_43 ? $signed(_spriteXRegs_43_T_2) : $signed({{16{_GEN_72[10]}},_GEN_72}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_451 = $signed(spriteXRegs_43) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_450); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_452 = $signed(spriteXRegs_43) >= 11'sh280 ? $signed(_spriteYRegs_43_T_2) : $signed(_GEN_73); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_453 = $signed(spriteXRegs_43) >= 11'sh280 ? lfsr_io_out_17[0] : _GEN_403; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _spriteYRegs_44_T_2 = 10'h64 + lfsr_io_out_28; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_1013 = {{16{spriteXRegs_44[10]}},spriteXRegs_44}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_44_T_2 = $signed(_GEN_1013) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_455 = spriteVisibleRegs_44 ? $signed(_spriteXRegs_44_T_2) : $signed({{16{_GEN_74[10]}},_GEN_74}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_456 = $signed(spriteXRegs_44) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_455); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_457 = $signed(spriteXRegs_44) >= 11'sh280 ? $signed(_spriteYRegs_44_T_2) : $signed(_GEN_75); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_458 = $signed(spriteXRegs_44) >= 11'sh280 ? lfsr_io_out_18[0] : _GEN_408; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _spriteYRegs_45_T_2 = 10'h64 + lfsr_io_out_29; // @[\\src\\main\\scala\\GameLogic.scala 423:63]
  wire [26:0] _GEN_1069 = {{16{spriteXRegs_45[10]}},spriteXRegs_45}; // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _spriteXRegs_45_T_2 = $signed(_GEN_1069) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 429:46]
  wire [26:0] _GEN_460 = spriteVisibleRegs_45 ? $signed(_spriteXRegs_45_T_2) : $signed({{16{_GEN_76[10]}},_GEN_76}); // @[\\src\\main\\scala\\GameLogic.scala 428:44 429:28]
  wire [26:0] _GEN_461 = $signed(spriteXRegs_45) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_460); // @[\\src\\main\\scala\\GameLogic.scala 421:41 422:28]
  wire [9:0] _GEN_462 = $signed(spriteXRegs_45) >= 11'sh280 ? $signed(_spriteYRegs_45_T_2) : $signed(_GEN_77); // @[\\src\\main\\scala\\GameLogic.scala 421:41 423:28]
  wire  _GEN_463 = $signed(spriteXRegs_45) >= 11'sh280 ? lfsr_io_out_19[0] : _GEN_413; // @[\\src\\main\\scala\\GameLogic.scala 421:41 426:40]
  wire [9:0] _extraLifeCnt_T_1 = extraLifeCnt + 10'h1; // @[\\src\\main\\scala\\GameLogic.scala 449:40]
  wire [10:0] _GEN_465 = extraLifeCnt == 10'h258 ? $signed(-11'sh20) : $signed(_GEN_14); // @[\\src\\main\\scala\\GameLogic.scala 443:38 444:27]
  wire  _GEN_466 = extraLifeCnt == 10'h258 | spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 443:38 445:33 125:34]
  wire [9:0] _GEN_467 = extraLifeCnt == 10'h258 ? $signed(lfsr_io_out_0) : $signed(_GEN_15); // @[\\src\\main\\scala\\GameLogic.scala 443:38 446:27]
  wire [9:0] _GEN_468 = extraLifeCnt == 10'h258 ? 10'h0 : _extraLifeCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 443:38 447:24 449:24]
  wire [10:0] _spriteXRegs_13_T_2 = $signed(spriteXRegs_13) + 11'sh2; // @[\\src\\main\\scala\\GameLogic.scala 452:46]
  wire [10:0] _GEN_469 = spriteVisibleRegs_13 ? $signed(_spriteXRegs_13_T_2) : $signed(_GEN_465); // @[\\src\\main\\scala\\GameLogic.scala 451:37 452:27]
  wire  _GEN_470 = $signed(spriteXRegs_13) >= 11'sh280 ? 1'h0 : _GEN_466; // @[\\src\\main\\scala\\GameLogic.scala 454:40 455:33]
  wire [26:0] _GEN_471 = _T ? $signed(_GEN_316) : $signed({{16{_GEN_18[10]}},_GEN_18}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_474 = _T ? _GEN_319 : spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_476 = _T ? $signed(_GEN_321) : $signed({{16{_GEN_20[10]}},_GEN_20}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_479 = _T ? _GEN_324 : spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_481 = _T ? $signed(_GEN_326) : $signed({{16{_GEN_22[10]}},_GEN_22}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_484 = _T ? _GEN_329 : spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_486 = _T ? $signed(_GEN_331) : $signed({{16{_GEN_24[10]}},_GEN_24}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_489 = _T ? _GEN_334 : spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_491 = _T ? $signed(_GEN_336) : $signed({{16{_GEN_26[10]}},_GEN_26}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_494 = _T ? _GEN_339 : spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_496 = _T ? $signed(_GEN_341) : $signed({{16{_GEN_28[10]}},_GEN_28}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_499 = _T ? _GEN_344 : spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_501 = _T ? $signed(_GEN_346) : $signed({{16{_GEN_30[10]}},_GEN_30}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_504 = _T ? _GEN_349 : spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_506 = _T ? $signed(_GEN_351) : $signed({{16{_GEN_32[10]}},_GEN_32}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_509 = _T ? _GEN_354 : spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_511 = _T ? $signed(_GEN_356) : $signed({{16{_GEN_34[10]}},_GEN_34}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_514 = _T ? _GEN_359 : spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_516 = _T ? $signed(_GEN_361) : $signed({{16{_GEN_36[10]}},_GEN_36}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_519 = _T ? _GEN_364 : spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 369:29 195:35]
  wire [26:0] _GEN_521 = _T ? $signed(_GEN_366) : $signed({{16{_GEN_38[10]}},_GEN_38}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_525 = _T ? $signed(_GEN_371) : $signed({{16{_GEN_40[10]}},_GEN_40}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_529 = _T ? $signed(_GEN_376) : $signed({{16{_GEN_42[10]}},_GEN_42}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_533 = _T ? $signed(_GEN_381) : $signed({{16{_GEN_44[10]}},_GEN_44}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_537 = _T ? $signed(_GEN_386) : $signed({{16{_GEN_46[10]}},_GEN_46}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_541 = _T ? $signed(_GEN_391) : $signed({{16{_GEN_48[10]}},_GEN_48}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_545 = _T ? $signed(_GEN_396) : $signed({{16{_GEN_50[10]}},_GEN_50}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_549 = _T ? $signed(_GEN_401) : $signed({{16{_GEN_52[10]}},_GEN_52}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_553 = _T ? $signed(_GEN_406) : $signed({{16{_GEN_54[10]}},_GEN_54}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_557 = _T ? $signed(_GEN_411) : $signed({{16{_GEN_56[10]}},_GEN_56}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_561 = _T ? $signed(_GEN_416) : $signed({{16{_GEN_58[10]}},_GEN_58}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_565 = _T ? $signed(_GEN_421) : $signed({{16{_GEN_60[10]}},_GEN_60}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_569 = _T ? $signed(_GEN_426) : $signed({{16{_GEN_62[10]}},_GEN_62}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_573 = _T ? $signed(_GEN_431) : $signed({{16{_GEN_64[10]}},_GEN_64}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_577 = _T ? $signed(_GEN_436) : $signed({{16{_GEN_66[10]}},_GEN_66}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_581 = _T ? $signed(_GEN_441) : $signed({{16{_GEN_68[10]}},_GEN_68}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_585 = _T ? $signed(_GEN_446) : $signed({{16{_GEN_70[10]}},_GEN_70}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_589 = _T ? $signed(_GEN_451) : $signed({{16{_GEN_72[10]}},_GEN_72}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_593 = _T ? $signed(_GEN_456) : $signed({{16{_GEN_74[10]}},_GEN_74}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire [26:0] _GEN_597 = _T ? $signed(_GEN_461) : $signed({{16{_GEN_76[10]}},_GEN_76}); // @[\\src\\main\\scala\\GameLogic.scala 369:29]
  wire  _GEN_602 = _T ? _GEN_470 : spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 369:29 125:34]
  wire  _T_69 = lvlReg == 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 460:19]
  wire  _T_72 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha; // @[\\src\\main\\scala\\GameLogic.scala 462:40]
  wire [5:0] _T_74 = 6'h10 + nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 463:34]
  wire  _GEN_608 = 6'h3 == _T_74 | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_609 = 6'h4 == _T_74 | spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_610 = 6'h5 == _T_74 | spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_611 = 6'h6 == _T_74 | spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_612 = 6'h7 == _T_74 | spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_613 = 6'h8 == _T_74 | spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_614 = 6'h9 == _T_74 | spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_615 = 6'ha == _T_74 | spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_616 = 6'hb == _T_74 | spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_617 = 6'hc == _T_74 | spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_618 = 6'hd == _T_74 | _GEN_602; // @[\\src\\main\\scala\\GameLogic.scala 463:{55,55}]
  wire  _GEN_619 = 6'he == _T_74 | spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_620 = 6'hf == _T_74 | spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_621 = 6'h10 == _T_74 | spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_622 = 6'h11 == _T_74 | spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_623 = 6'h12 == _T_74 | spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_624 = 6'h13 == _T_74 | spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_625 = 6'h14 == _T_74 | spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_626 = 6'h15 == _T_74 | spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_627 = 6'h16 == _T_74 | spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_628 = 6'h17 == _T_74 | spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_629 = 6'h18 == _T_74 | spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_630 = 6'h19 == _T_74 | spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_631 = 6'h1a == _T_74 | spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_632 = 6'h1b == _T_74 | spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_633 = 6'h1c == _T_74 | spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_634 = 6'h1d == _T_74 | spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_635 = 6'h1e == _T_74 | spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_636 = 6'h1f == _T_74 | spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_637 = 6'h20 == _T_74 | spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_638 = 6'h21 == _T_74 | spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_639 = 6'h22 == _T_74 | spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_640 = 6'h23 == _T_74 | spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_641 = 6'h24 == _T_74 | spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_642 = 6'h25 == _T_74 | spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_643 = 6'h26 == _T_74 | spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_644 = 6'h27 == _T_74 | spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_645 = 6'h28 == _T_74 | spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_646 = 6'h29 == _T_74 | spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_647 = 6'h2a == _T_74 | spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_648 = 6'h2b == _T_74 | spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_649 = 6'h2c == _T_74 | spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_650 = 6'h2d == _T_74 | spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_651 = 6'h2e == _T_74 | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_652 = 6'h2f == _T_74 | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_653 = 6'h30 == _T_74 | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_654 = 6'h31 == _T_74 | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_655 = 6'h32 == _T_74 | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_656 = 6'h33 == _T_74 | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_657 = 6'h34 == _T_74 | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_658 = 6'h35 == _T_74 | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_659 = 6'h36 == _T_74 | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_660 = 6'h37 == _T_74 | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_661 = 6'h38 == _T_74 | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_662 = 6'h39 == _T_74 | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_666 = 6'h3d == _T_74 | _GEN_195; // @[\\src\\main\\scala\\GameLogic.scala 463:{55,55}]
  wire  _GEN_667 = 6'h3e == _T_74 | _GEN_196; // @[\\src\\main\\scala\\GameLogic.scala 463:{55,55}]
  wire  _GEN_668 = 6'h3f == _T_74 | _GEN_197; // @[\\src\\main\\scala\\GameLogic.scala 463:{55,55}]
  wire [6:0] _GEN_2383 = {{1'd0}, _T_74}; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_669 = 7'h40 == _GEN_2383 | spriteVisibleRegs_64; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_670 = 7'h41 == _GEN_2383 | spriteVisibleRegs_65; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_671 = 7'h42 == _GEN_2383 | spriteVisibleRegs_66; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_672 = 7'h43 == _GEN_2383 | spriteVisibleRegs_67; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_673 = 7'h44 == _GEN_2383 | spriteVisibleRegs_68; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_674 = 7'h45 == _GEN_2383 | spriteVisibleRegs_69; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_675 = 7'h46 == _GEN_2383 | spriteVisibleRegs_70; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_676 = 7'h47 == _GEN_2383 | spriteVisibleRegs_71; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_677 = 7'h48 == _GEN_2383 | spriteVisibleRegs_72; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_678 = 7'h49 == _GEN_2383 | spriteVisibleRegs_73; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_679 = 7'h4a == _GEN_2383 | spriteVisibleRegs_74; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_680 = 7'h4b == _GEN_2383 | spriteVisibleRegs_75; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_681 = 7'h4c == _GEN_2383 | spriteVisibleRegs_76; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_682 = 7'h4d == _GEN_2383 | spriteVisibleRegs_77; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_683 = 7'h4e == _GEN_2383 | spriteVisibleRegs_78; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_684 = 7'h4f == _GEN_2383 | spriteVisibleRegs_79; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_685 = 7'h50 == _GEN_2383 | spriteVisibleRegs_80; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_686 = 7'h51 == _GEN_2383 | spriteVisibleRegs_81; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_687 = 7'h52 == _GEN_2383 | spriteVisibleRegs_82; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_688 = 7'h53 == _GEN_2383 | spriteVisibleRegs_83; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_689 = 7'h54 == _GEN_2383 | spriteVisibleRegs_84; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_690 = 7'h55 == _GEN_2383 | spriteVisibleRegs_85; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_691 = 7'h56 == _GEN_2383 | spriteVisibleRegs_86; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_692 = 7'h57 == _GEN_2383 | spriteVisibleRegs_87; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_693 = 7'h58 == _GEN_2383 | spriteVisibleRegs_88; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_694 = 7'h59 == _GEN_2383 | spriteVisibleRegs_89; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_695 = 7'h5a == _GEN_2383 | spriteVisibleRegs_90; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_696 = 7'h5b == _GEN_2383 | spriteVisibleRegs_91; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_697 = 7'h5c == _GEN_2383 | spriteVisibleRegs_92; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_698 = 7'h5d == _GEN_2383 | spriteVisibleRegs_93; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_699 = 7'h5e == _GEN_2383 | spriteVisibleRegs_94; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_700 = 7'h5f == _GEN_2383 | spriteVisibleRegs_95; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_701 = 7'h60 == _GEN_2383 | spriteVisibleRegs_96; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_702 = 7'h61 == _GEN_2383 | spriteVisibleRegs_97; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_703 = 7'h62 == _GEN_2383 | spriteVisibleRegs_98; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire  _GEN_704 = 7'h63 == _GEN_2383 | spriteVisibleRegs_99; // @[\\src\\main\\scala\\GameLogic.scala 125:34 463:{55,55}]
  wire [5:0] _nextSpriteToSpawn_T_1 = nextSpriteToSpawn + 6'h1; // @[\\src\\main\\scala\\GameLogic.scala 464:50]
  wire [7:0] _spawnDelayCounter_T_1 = spawnDelayCounter - 8'h1; // @[\\src\\main\\scala\\GameLogic.scala 467:50]
  wire [7:0] _GEN_705 = spawnDelayCounter > 8'h0 ? _spawnDelayCounter_T_1 : spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 466:45 467:29 243:34]
  wire  _GEN_709 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_608 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_710 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_609 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_711 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_610 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_712 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_611 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_713 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_612 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_714 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_613 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_715 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_614 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_716 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_615 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_717 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_616 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_718 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_617 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_719 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_618 : _GEN_602; // @[\\src\\main\\scala\\GameLogic.scala 462:69]
  wire  _GEN_720 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_619 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_721 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_620 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_722 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_621 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_723 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_622 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_724 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_623 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_725 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_624 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_726 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_625 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_727 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_626 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_728 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_627 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_729 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_628 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_730 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_629 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_731 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_630 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_732 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_631 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_733 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_632 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_734 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_633 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_735 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_634 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_736 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_635 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_737 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_636 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_738 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_637 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_739 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_638 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_740 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_639 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_741 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_640 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_742 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_641 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_743 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_642 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_744 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_643 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_745 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_644 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_746 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_645 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_747 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_646 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_748 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_647 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_749 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_648 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_750 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_649 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_751 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_650 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_752 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_651 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_753 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_652 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_754 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_653 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_755 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_654 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_756 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_655 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_757 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_656 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_758 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_657 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_759 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_658 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_760 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_659 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_761 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_660 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_762 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_661 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_763 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_662 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_767 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_666 : _GEN_195; // @[\\src\\main\\scala\\GameLogic.scala 462:69]
  wire  _GEN_768 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_667 : _GEN_196; // @[\\src\\main\\scala\\GameLogic.scala 462:69]
  wire  _GEN_769 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_668 : _GEN_197; // @[\\src\\main\\scala\\GameLogic.scala 462:69]
  wire  _GEN_770 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_669 : spriteVisibleRegs_64; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_771 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_670 : spriteVisibleRegs_65; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_772 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_671 : spriteVisibleRegs_66; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_773 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_672 : spriteVisibleRegs_67; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_774 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_673 : spriteVisibleRegs_68; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_775 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_674 : spriteVisibleRegs_69; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_776 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_675 : spriteVisibleRegs_70; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_777 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_676 : spriteVisibleRegs_71; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_778 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_677 : spriteVisibleRegs_72; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_779 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_678 : spriteVisibleRegs_73; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_780 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_679 : spriteVisibleRegs_74; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_781 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_680 : spriteVisibleRegs_75; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_782 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_681 : spriteVisibleRegs_76; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_783 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_682 : spriteVisibleRegs_77; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_784 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_683 : spriteVisibleRegs_78; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_785 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_684 : spriteVisibleRegs_79; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_786 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_685 : spriteVisibleRegs_80; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_787 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_686 : spriteVisibleRegs_81; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_788 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_687 : spriteVisibleRegs_82; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_789 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_688 : spriteVisibleRegs_83; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_790 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_689 : spriteVisibleRegs_84; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_791 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_690 : spriteVisibleRegs_85; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_792 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_691 : spriteVisibleRegs_86; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_793 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_692 : spriteVisibleRegs_87; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_794 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_693 : spriteVisibleRegs_88; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_795 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_694 : spriteVisibleRegs_89; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_796 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_695 : spriteVisibleRegs_90; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_797 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_696 : spriteVisibleRegs_91; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_798 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_697 : spriteVisibleRegs_92; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_799 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_698 : spriteVisibleRegs_93; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_800 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_699 : spriteVisibleRegs_94; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_801 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_700 : spriteVisibleRegs_95; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_802 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_701 : spriteVisibleRegs_96; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_803 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_702 : spriteVisibleRegs_97; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_804 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_703 : spriteVisibleRegs_98; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire  _GEN_805 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_704 : spriteVisibleRegs_99; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:69]
  wire [5:0] _GEN_806 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _nextSpriteToSpawn_T_1 :
    nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 462:69 464:29 244:34]
  wire [7:0] _GEN_807 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? 8'h1e : _GEN_705; // @[\\src\\main\\scala\\GameLogic.scala 462:69 465:29]
  wire  _T_76 = lvlReg == 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 469:25]
  wire [5:0] _T_81 = 6'h1a + nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 472:34]
  wire  _GEN_811 = 6'h3 == _T_81 | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_812 = 6'h4 == _T_81 | spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_813 = 6'h5 == _T_81 | spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_814 = 6'h6 == _T_81 | spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_815 = 6'h7 == _T_81 | spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_816 = 6'h8 == _T_81 | spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_817 = 6'h9 == _T_81 | spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_818 = 6'ha == _T_81 | spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_819 = 6'hb == _T_81 | spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_820 = 6'hc == _T_81 | spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_821 = 6'hd == _T_81 | _GEN_602; // @[\\src\\main\\scala\\GameLogic.scala 472:{55,55}]
  wire  _GEN_822 = 6'he == _T_81 | spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_823 = 6'hf == _T_81 | spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_824 = 6'h10 == _T_81 | spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_825 = 6'h11 == _T_81 | spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_826 = 6'h12 == _T_81 | spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_827 = 6'h13 == _T_81 | spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_828 = 6'h14 == _T_81 | spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_829 = 6'h15 == _T_81 | spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_830 = 6'h16 == _T_81 | spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_831 = 6'h17 == _T_81 | spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_832 = 6'h18 == _T_81 | spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_833 = 6'h19 == _T_81 | spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_834 = 6'h1a == _T_81 | spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_835 = 6'h1b == _T_81 | spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_836 = 6'h1c == _T_81 | spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_837 = 6'h1d == _T_81 | spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_838 = 6'h1e == _T_81 | spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_839 = 6'h1f == _T_81 | spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_840 = 6'h20 == _T_81 | spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_841 = 6'h21 == _T_81 | spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_842 = 6'h22 == _T_81 | spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_843 = 6'h23 == _T_81 | spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_844 = 6'h24 == _T_81 | spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_845 = 6'h25 == _T_81 | spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_846 = 6'h26 == _T_81 | spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_847 = 6'h27 == _T_81 | spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_848 = 6'h28 == _T_81 | spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_849 = 6'h29 == _T_81 | spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_850 = 6'h2a == _T_81 | spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_851 = 6'h2b == _T_81 | spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_852 = 6'h2c == _T_81 | spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_853 = 6'h2d == _T_81 | spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_854 = 6'h2e == _T_81 | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_855 = 6'h2f == _T_81 | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_856 = 6'h30 == _T_81 | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_857 = 6'h31 == _T_81 | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_858 = 6'h32 == _T_81 | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_859 = 6'h33 == _T_81 | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_860 = 6'h34 == _T_81 | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_861 = 6'h35 == _T_81 | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_862 = 6'h36 == _T_81 | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_863 = 6'h37 == _T_81 | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_864 = 6'h38 == _T_81 | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_865 = 6'h39 == _T_81 | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_869 = 6'h3d == _T_81 | _GEN_195; // @[\\src\\main\\scala\\GameLogic.scala 472:{55,55}]
  wire  _GEN_870 = 6'h3e == _T_81 | _GEN_196; // @[\\src\\main\\scala\\GameLogic.scala 472:{55,55}]
  wire  _GEN_871 = 6'h3f == _T_81 | _GEN_197; // @[\\src\\main\\scala\\GameLogic.scala 472:{55,55}]
  wire [6:0] _GEN_2513 = {{1'd0}, _T_81}; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_872 = 7'h40 == _GEN_2513 | spriteVisibleRegs_64; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_873 = 7'h41 == _GEN_2513 | spriteVisibleRegs_65; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_874 = 7'h42 == _GEN_2513 | spriteVisibleRegs_66; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_875 = 7'h43 == _GEN_2513 | spriteVisibleRegs_67; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_876 = 7'h44 == _GEN_2513 | spriteVisibleRegs_68; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_877 = 7'h45 == _GEN_2513 | spriteVisibleRegs_69; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_878 = 7'h46 == _GEN_2513 | spriteVisibleRegs_70; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_879 = 7'h47 == _GEN_2513 | spriteVisibleRegs_71; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_880 = 7'h48 == _GEN_2513 | spriteVisibleRegs_72; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_881 = 7'h49 == _GEN_2513 | spriteVisibleRegs_73; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_882 = 7'h4a == _GEN_2513 | spriteVisibleRegs_74; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_883 = 7'h4b == _GEN_2513 | spriteVisibleRegs_75; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_884 = 7'h4c == _GEN_2513 | spriteVisibleRegs_76; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_885 = 7'h4d == _GEN_2513 | spriteVisibleRegs_77; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_886 = 7'h4e == _GEN_2513 | spriteVisibleRegs_78; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_887 = 7'h4f == _GEN_2513 | spriteVisibleRegs_79; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_888 = 7'h50 == _GEN_2513 | spriteVisibleRegs_80; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_889 = 7'h51 == _GEN_2513 | spriteVisibleRegs_81; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_890 = 7'h52 == _GEN_2513 | spriteVisibleRegs_82; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_891 = 7'h53 == _GEN_2513 | spriteVisibleRegs_83; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_892 = 7'h54 == _GEN_2513 | spriteVisibleRegs_84; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_893 = 7'h55 == _GEN_2513 | spriteVisibleRegs_85; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_894 = 7'h56 == _GEN_2513 | spriteVisibleRegs_86; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_895 = 7'h57 == _GEN_2513 | spriteVisibleRegs_87; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_896 = 7'h58 == _GEN_2513 | spriteVisibleRegs_88; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_897 = 7'h59 == _GEN_2513 | spriteVisibleRegs_89; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_898 = 7'h5a == _GEN_2513 | spriteVisibleRegs_90; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_899 = 7'h5b == _GEN_2513 | spriteVisibleRegs_91; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_900 = 7'h5c == _GEN_2513 | spriteVisibleRegs_92; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_901 = 7'h5d == _GEN_2513 | spriteVisibleRegs_93; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_902 = 7'h5e == _GEN_2513 | spriteVisibleRegs_94; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_903 = 7'h5f == _GEN_2513 | spriteVisibleRegs_95; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_904 = 7'h60 == _GEN_2513 | spriteVisibleRegs_96; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_905 = 7'h61 == _GEN_2513 | spriteVisibleRegs_97; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_906 = 7'h62 == _GEN_2513 | spriteVisibleRegs_98; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_907 = 7'h63 == _GEN_2513 | spriteVisibleRegs_99; // @[\\src\\main\\scala\\GameLogic.scala 125:34 472:{55,55}]
  wire  _GEN_912 = _T_72 ? _GEN_811 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_913 = _T_72 ? _GEN_812 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_914 = _T_72 ? _GEN_813 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_915 = _T_72 ? _GEN_814 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_916 = _T_72 ? _GEN_815 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_917 = _T_72 ? _GEN_816 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_918 = _T_72 ? _GEN_817 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_919 = _T_72 ? _GEN_818 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_920 = _T_72 ? _GEN_819 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_921 = _T_72 ? _GEN_820 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_922 = _T_72 ? _GEN_821 : _GEN_602; // @[\\src\\main\\scala\\GameLogic.scala 471:69]
  wire  _GEN_923 = _T_72 ? _GEN_822 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_924 = _T_72 ? _GEN_823 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_925 = _T_72 ? _GEN_824 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_926 = _T_72 ? _GEN_825 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_927 = _T_72 ? _GEN_826 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_928 = _T_72 ? _GEN_827 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_929 = _T_72 ? _GEN_828 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_930 = _T_72 ? _GEN_829 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_931 = _T_72 ? _GEN_830 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_932 = _T_72 ? _GEN_831 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_933 = _T_72 ? _GEN_832 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_934 = _T_72 ? _GEN_833 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_935 = _T_72 ? _GEN_834 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_936 = _T_72 ? _GEN_835 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_937 = _T_72 ? _GEN_836 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_938 = _T_72 ? _GEN_837 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_939 = _T_72 ? _GEN_838 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_940 = _T_72 ? _GEN_839 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_941 = _T_72 ? _GEN_840 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_942 = _T_72 ? _GEN_841 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_943 = _T_72 ? _GEN_842 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_944 = _T_72 ? _GEN_843 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_945 = _T_72 ? _GEN_844 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_946 = _T_72 ? _GEN_845 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_947 = _T_72 ? _GEN_846 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_948 = _T_72 ? _GEN_847 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_949 = _T_72 ? _GEN_848 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_950 = _T_72 ? _GEN_849 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_951 = _T_72 ? _GEN_850 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_952 = _T_72 ? _GEN_851 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_953 = _T_72 ? _GEN_852 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_954 = _T_72 ? _GEN_853 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_955 = _T_72 ? _GEN_854 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_956 = _T_72 ? _GEN_855 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_957 = _T_72 ? _GEN_856 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_958 = _T_72 ? _GEN_857 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_959 = _T_72 ? _GEN_858 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_960 = _T_72 ? _GEN_859 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_961 = _T_72 ? _GEN_860 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_962 = _T_72 ? _GEN_861 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_963 = _T_72 ? _GEN_862 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_964 = _T_72 ? _GEN_863 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_965 = _T_72 ? _GEN_864 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_966 = _T_72 ? _GEN_865 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_970 = _T_72 ? _GEN_869 : _GEN_195; // @[\\src\\main\\scala\\GameLogic.scala 471:69]
  wire  _GEN_971 = _T_72 ? _GEN_870 : _GEN_196; // @[\\src\\main\\scala\\GameLogic.scala 471:69]
  wire  _GEN_972 = _T_72 ? _GEN_871 : _GEN_197; // @[\\src\\main\\scala\\GameLogic.scala 471:69]
  wire  _GEN_973 = _T_72 ? _GEN_872 : spriteVisibleRegs_64; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_974 = _T_72 ? _GEN_873 : spriteVisibleRegs_65; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_975 = _T_72 ? _GEN_874 : spriteVisibleRegs_66; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_976 = _T_72 ? _GEN_875 : spriteVisibleRegs_67; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_977 = _T_72 ? _GEN_876 : spriteVisibleRegs_68; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_978 = _T_72 ? _GEN_877 : spriteVisibleRegs_69; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_979 = _T_72 ? _GEN_878 : spriteVisibleRegs_70; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_980 = _T_72 ? _GEN_879 : spriteVisibleRegs_71; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_981 = _T_72 ? _GEN_880 : spriteVisibleRegs_72; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_982 = _T_72 ? _GEN_881 : spriteVisibleRegs_73; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_983 = _T_72 ? _GEN_882 : spriteVisibleRegs_74; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_984 = _T_72 ? _GEN_883 : spriteVisibleRegs_75; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_985 = _T_72 ? _GEN_884 : spriteVisibleRegs_76; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_986 = _T_72 ? _GEN_885 : spriteVisibleRegs_77; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_987 = _T_72 ? _GEN_886 : spriteVisibleRegs_78; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_988 = _T_72 ? _GEN_887 : spriteVisibleRegs_79; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_989 = _T_72 ? _GEN_888 : spriteVisibleRegs_80; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_990 = _T_72 ? _GEN_889 : spriteVisibleRegs_81; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_991 = _T_72 ? _GEN_890 : spriteVisibleRegs_82; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_992 = _T_72 ? _GEN_891 : spriteVisibleRegs_83; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_993 = _T_72 ? _GEN_892 : spriteVisibleRegs_84; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_994 = _T_72 ? _GEN_893 : spriteVisibleRegs_85; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_995 = _T_72 ? _GEN_894 : spriteVisibleRegs_86; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_996 = _T_72 ? _GEN_895 : spriteVisibleRegs_87; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_997 = _T_72 ? _GEN_896 : spriteVisibleRegs_88; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_998 = _T_72 ? _GEN_897 : spriteVisibleRegs_89; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_999 = _T_72 ? _GEN_898 : spriteVisibleRegs_90; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_1000 = _T_72 ? _GEN_899 : spriteVisibleRegs_91; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_1001 = _T_72 ? _GEN_900 : spriteVisibleRegs_92; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_1002 = _T_72 ? _GEN_901 : spriteVisibleRegs_93; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_1003 = _T_72 ? _GEN_902 : spriteVisibleRegs_94; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_1004 = _T_72 ? _GEN_903 : spriteVisibleRegs_95; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_1005 = _T_72 ? _GEN_904 : spriteVisibleRegs_96; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_1006 = _T_72 ? _GEN_905 : spriteVisibleRegs_97; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_1007 = _T_72 ? _GEN_906 : spriteVisibleRegs_98; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire  _GEN_1008 = _T_72 ? _GEN_907 : spriteVisibleRegs_99; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:69]
  wire [7:0] _GEN_1010 = _T_72 ? 8'h19 : _GEN_705; // @[\\src\\main\\scala\\GameLogic.scala 471:69 474:29]
  wire  _T_83 = lvlReg == 2'h3; // @[\\src\\main\\scala\\GameLogic.scala 478:25]
  wire [5:0] _T_88 = 6'h24 + nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 481:34]
  wire  _GEN_1014 = 6'h3 == _T_88 | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1015 = 6'h4 == _T_88 | spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1016 = 6'h5 == _T_88 | spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1017 = 6'h6 == _T_88 | spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1018 = 6'h7 == _T_88 | spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1019 = 6'h8 == _T_88 | spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1020 = 6'h9 == _T_88 | spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1021 = 6'ha == _T_88 | spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1022 = 6'hb == _T_88 | spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1023 = 6'hc == _T_88 | spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1024 = 6'hd == _T_88 | _GEN_602; // @[\\src\\main\\scala\\GameLogic.scala 481:{55,55}]
  wire  _GEN_1025 = 6'he == _T_88 | spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1026 = 6'hf == _T_88 | spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1027 = 6'h10 == _T_88 | spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1028 = 6'h11 == _T_88 | spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1029 = 6'h12 == _T_88 | spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1030 = 6'h13 == _T_88 | spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1031 = 6'h14 == _T_88 | spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1032 = 6'h15 == _T_88 | spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1033 = 6'h16 == _T_88 | spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1034 = 6'h17 == _T_88 | spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1035 = 6'h18 == _T_88 | spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1036 = 6'h19 == _T_88 | spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1037 = 6'h1a == _T_88 | spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1038 = 6'h1b == _T_88 | spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1039 = 6'h1c == _T_88 | spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1040 = 6'h1d == _T_88 | spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1041 = 6'h1e == _T_88 | spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1042 = 6'h1f == _T_88 | spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1043 = 6'h20 == _T_88 | spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1044 = 6'h21 == _T_88 | spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1045 = 6'h22 == _T_88 | spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1046 = 6'h23 == _T_88 | spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1047 = 6'h24 == _T_88 | spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1048 = 6'h25 == _T_88 | spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1049 = 6'h26 == _T_88 | spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1050 = 6'h27 == _T_88 | spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1051 = 6'h28 == _T_88 | spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1052 = 6'h29 == _T_88 | spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1053 = 6'h2a == _T_88 | spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1054 = 6'h2b == _T_88 | spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1055 = 6'h2c == _T_88 | spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1056 = 6'h2d == _T_88 | spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1057 = 6'h2e == _T_88 | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1058 = 6'h2f == _T_88 | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1059 = 6'h30 == _T_88 | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1060 = 6'h31 == _T_88 | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1061 = 6'h32 == _T_88 | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1062 = 6'h33 == _T_88 | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1063 = 6'h34 == _T_88 | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1064 = 6'h35 == _T_88 | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1065 = 6'h36 == _T_88 | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1066 = 6'h37 == _T_88 | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1067 = 6'h38 == _T_88 | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1068 = 6'h39 == _T_88 | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1072 = 6'h3d == _T_88 | _GEN_195; // @[\\src\\main\\scala\\GameLogic.scala 481:{55,55}]
  wire  _GEN_1073 = 6'h3e == _T_88 | _GEN_196; // @[\\src\\main\\scala\\GameLogic.scala 481:{55,55}]
  wire  _GEN_1074 = 6'h3f == _T_88 | _GEN_197; // @[\\src\\main\\scala\\GameLogic.scala 481:{55,55}]
  wire [6:0] _GEN_2643 = {{1'd0}, _T_88}; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1075 = 7'h40 == _GEN_2643 | spriteVisibleRegs_64; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1076 = 7'h41 == _GEN_2643 | spriteVisibleRegs_65; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1077 = 7'h42 == _GEN_2643 | spriteVisibleRegs_66; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1078 = 7'h43 == _GEN_2643 | spriteVisibleRegs_67; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1079 = 7'h44 == _GEN_2643 | spriteVisibleRegs_68; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1080 = 7'h45 == _GEN_2643 | spriteVisibleRegs_69; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1081 = 7'h46 == _GEN_2643 | spriteVisibleRegs_70; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1082 = 7'h47 == _GEN_2643 | spriteVisibleRegs_71; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1083 = 7'h48 == _GEN_2643 | spriteVisibleRegs_72; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1084 = 7'h49 == _GEN_2643 | spriteVisibleRegs_73; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1085 = 7'h4a == _GEN_2643 | spriteVisibleRegs_74; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1086 = 7'h4b == _GEN_2643 | spriteVisibleRegs_75; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1087 = 7'h4c == _GEN_2643 | spriteVisibleRegs_76; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1088 = 7'h4d == _GEN_2643 | spriteVisibleRegs_77; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1089 = 7'h4e == _GEN_2643 | spriteVisibleRegs_78; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1090 = 7'h4f == _GEN_2643 | spriteVisibleRegs_79; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1091 = 7'h50 == _GEN_2643 | spriteVisibleRegs_80; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1092 = 7'h51 == _GEN_2643 | spriteVisibleRegs_81; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1093 = 7'h52 == _GEN_2643 | spriteVisibleRegs_82; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1094 = 7'h53 == _GEN_2643 | spriteVisibleRegs_83; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1095 = 7'h54 == _GEN_2643 | spriteVisibleRegs_84; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1096 = 7'h55 == _GEN_2643 | spriteVisibleRegs_85; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1097 = 7'h56 == _GEN_2643 | spriteVisibleRegs_86; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1098 = 7'h57 == _GEN_2643 | spriteVisibleRegs_87; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1099 = 7'h58 == _GEN_2643 | spriteVisibleRegs_88; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1100 = 7'h59 == _GEN_2643 | spriteVisibleRegs_89; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1101 = 7'h5a == _GEN_2643 | spriteVisibleRegs_90; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1102 = 7'h5b == _GEN_2643 | spriteVisibleRegs_91; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1103 = 7'h5c == _GEN_2643 | spriteVisibleRegs_92; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1104 = 7'h5d == _GEN_2643 | spriteVisibleRegs_93; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1105 = 7'h5e == _GEN_2643 | spriteVisibleRegs_94; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1106 = 7'h5f == _GEN_2643 | spriteVisibleRegs_95; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1107 = 7'h60 == _GEN_2643 | spriteVisibleRegs_96; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1108 = 7'h61 == _GEN_2643 | spriteVisibleRegs_97; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1109 = 7'h62 == _GEN_2643 | spriteVisibleRegs_98; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1110 = 7'h63 == _GEN_2643 | spriteVisibleRegs_99; // @[\\src\\main\\scala\\GameLogic.scala 125:34 481:{55,55}]
  wire  _GEN_1115 = _T_72 ? _GEN_1014 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1116 = _T_72 ? _GEN_1015 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1117 = _T_72 ? _GEN_1016 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1118 = _T_72 ? _GEN_1017 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1119 = _T_72 ? _GEN_1018 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1120 = _T_72 ? _GEN_1019 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1121 = _T_72 ? _GEN_1020 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1122 = _T_72 ? _GEN_1021 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1123 = _T_72 ? _GEN_1022 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1124 = _T_72 ? _GEN_1023 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1125 = _T_72 ? _GEN_1024 : _GEN_602; // @[\\src\\main\\scala\\GameLogic.scala 480:69]
  wire  _GEN_1126 = _T_72 ? _GEN_1025 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1127 = _T_72 ? _GEN_1026 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1128 = _T_72 ? _GEN_1027 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1129 = _T_72 ? _GEN_1028 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1130 = _T_72 ? _GEN_1029 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1131 = _T_72 ? _GEN_1030 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1132 = _T_72 ? _GEN_1031 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1133 = _T_72 ? _GEN_1032 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1134 = _T_72 ? _GEN_1033 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1135 = _T_72 ? _GEN_1034 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1136 = _T_72 ? _GEN_1035 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1137 = _T_72 ? _GEN_1036 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1138 = _T_72 ? _GEN_1037 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1139 = _T_72 ? _GEN_1038 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1140 = _T_72 ? _GEN_1039 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1141 = _T_72 ? _GEN_1040 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1142 = _T_72 ? _GEN_1041 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1143 = _T_72 ? _GEN_1042 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1144 = _T_72 ? _GEN_1043 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1145 = _T_72 ? _GEN_1044 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1146 = _T_72 ? _GEN_1045 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1147 = _T_72 ? _GEN_1046 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1148 = _T_72 ? _GEN_1047 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1149 = _T_72 ? _GEN_1048 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1150 = _T_72 ? _GEN_1049 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1151 = _T_72 ? _GEN_1050 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1152 = _T_72 ? _GEN_1051 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1153 = _T_72 ? _GEN_1052 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1154 = _T_72 ? _GEN_1053 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1155 = _T_72 ? _GEN_1054 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1156 = _T_72 ? _GEN_1055 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1157 = _T_72 ? _GEN_1056 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1158 = _T_72 ? _GEN_1057 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1159 = _T_72 ? _GEN_1058 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1160 = _T_72 ? _GEN_1059 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1161 = _T_72 ? _GEN_1060 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1162 = _T_72 ? _GEN_1061 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1163 = _T_72 ? _GEN_1062 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1164 = _T_72 ? _GEN_1063 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1165 = _T_72 ? _GEN_1064 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1166 = _T_72 ? _GEN_1065 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1167 = _T_72 ? _GEN_1066 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1168 = _T_72 ? _GEN_1067 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1169 = _T_72 ? _GEN_1068 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1173 = _T_72 ? _GEN_1072 : _GEN_195; // @[\\src\\main\\scala\\GameLogic.scala 480:69]
  wire  _GEN_1174 = _T_72 ? _GEN_1073 : _GEN_196; // @[\\src\\main\\scala\\GameLogic.scala 480:69]
  wire  _GEN_1175 = _T_72 ? _GEN_1074 : _GEN_197; // @[\\src\\main\\scala\\GameLogic.scala 480:69]
  wire  _GEN_1176 = _T_72 ? _GEN_1075 : spriteVisibleRegs_64; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1177 = _T_72 ? _GEN_1076 : spriteVisibleRegs_65; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1178 = _T_72 ? _GEN_1077 : spriteVisibleRegs_66; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1179 = _T_72 ? _GEN_1078 : spriteVisibleRegs_67; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1180 = _T_72 ? _GEN_1079 : spriteVisibleRegs_68; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1181 = _T_72 ? _GEN_1080 : spriteVisibleRegs_69; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1182 = _T_72 ? _GEN_1081 : spriteVisibleRegs_70; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1183 = _T_72 ? _GEN_1082 : spriteVisibleRegs_71; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1184 = _T_72 ? _GEN_1083 : spriteVisibleRegs_72; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1185 = _T_72 ? _GEN_1084 : spriteVisibleRegs_73; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1186 = _T_72 ? _GEN_1085 : spriteVisibleRegs_74; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1187 = _T_72 ? _GEN_1086 : spriteVisibleRegs_75; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1188 = _T_72 ? _GEN_1087 : spriteVisibleRegs_76; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1189 = _T_72 ? _GEN_1088 : spriteVisibleRegs_77; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1190 = _T_72 ? _GEN_1089 : spriteVisibleRegs_78; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1191 = _T_72 ? _GEN_1090 : spriteVisibleRegs_79; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1192 = _T_72 ? _GEN_1091 : spriteVisibleRegs_80; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1193 = _T_72 ? _GEN_1092 : spriteVisibleRegs_81; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1194 = _T_72 ? _GEN_1093 : spriteVisibleRegs_82; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1195 = _T_72 ? _GEN_1094 : spriteVisibleRegs_83; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1196 = _T_72 ? _GEN_1095 : spriteVisibleRegs_84; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1197 = _T_72 ? _GEN_1096 : spriteVisibleRegs_85; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1198 = _T_72 ? _GEN_1097 : spriteVisibleRegs_86; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1199 = _T_72 ? _GEN_1098 : spriteVisibleRegs_87; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1200 = _T_72 ? _GEN_1099 : spriteVisibleRegs_88; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1201 = _T_72 ? _GEN_1100 : spriteVisibleRegs_89; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1202 = _T_72 ? _GEN_1101 : spriteVisibleRegs_90; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1203 = _T_72 ? _GEN_1102 : spriteVisibleRegs_91; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1204 = _T_72 ? _GEN_1103 : spriteVisibleRegs_92; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1205 = _T_72 ? _GEN_1104 : spriteVisibleRegs_93; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1206 = _T_72 ? _GEN_1105 : spriteVisibleRegs_94; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1207 = _T_72 ? _GEN_1106 : spriteVisibleRegs_95; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1208 = _T_72 ? _GEN_1107 : spriteVisibleRegs_96; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1209 = _T_72 ? _GEN_1108 : spriteVisibleRegs_97; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1210 = _T_72 ? _GEN_1109 : spriteVisibleRegs_98; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire  _GEN_1211 = _T_72 ? _GEN_1110 : spriteVisibleRegs_99; // @[\\src\\main\\scala\\GameLogic.scala 125:34 480:69]
  wire [7:0] _GEN_1213 = _T_72 ? 8'h14 : _GEN_705; // @[\\src\\main\\scala\\GameLogic.scala 480:69 483:29]
  wire  _GEN_1217 = lvlReg == 2'h3 ? _GEN_1115 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1218 = lvlReg == 2'h3 ? _GEN_1116 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1219 = lvlReg == 2'h3 ? _GEN_1117 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1220 = lvlReg == 2'h3 ? _GEN_1118 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1221 = lvlReg == 2'h3 ? _GEN_1119 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1222 = lvlReg == 2'h3 ? _GEN_1120 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1223 = lvlReg == 2'h3 ? _GEN_1121 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1224 = lvlReg == 2'h3 ? _GEN_1122 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1225 = lvlReg == 2'h3 ? _GEN_1123 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1226 = lvlReg == 2'h3 ? _GEN_1124 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1227 = lvlReg == 2'h3 ? _GEN_1125 : _GEN_602; // @[\\src\\main\\scala\\GameLogic.scala 478:34]
  wire  _GEN_1228 = lvlReg == 2'h3 ? _GEN_1126 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1229 = lvlReg == 2'h3 ? _GEN_1127 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1230 = lvlReg == 2'h3 ? _GEN_1128 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1231 = lvlReg == 2'h3 ? _GEN_1129 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1232 = lvlReg == 2'h3 ? _GEN_1130 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1233 = lvlReg == 2'h3 ? _GEN_1131 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1234 = lvlReg == 2'h3 ? _GEN_1132 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1235 = lvlReg == 2'h3 ? _GEN_1133 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1236 = lvlReg == 2'h3 ? _GEN_1134 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1237 = lvlReg == 2'h3 ? _GEN_1135 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1238 = lvlReg == 2'h3 ? _GEN_1136 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1239 = lvlReg == 2'h3 ? _GEN_1137 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1240 = lvlReg == 2'h3 ? _GEN_1138 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1241 = lvlReg == 2'h3 ? _GEN_1139 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1242 = lvlReg == 2'h3 ? _GEN_1140 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1243 = lvlReg == 2'h3 ? _GEN_1141 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1244 = lvlReg == 2'h3 ? _GEN_1142 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1245 = lvlReg == 2'h3 ? _GEN_1143 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1246 = lvlReg == 2'h3 ? _GEN_1144 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1247 = lvlReg == 2'h3 ? _GEN_1145 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1248 = lvlReg == 2'h3 ? _GEN_1146 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1249 = lvlReg == 2'h3 ? _GEN_1147 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1250 = lvlReg == 2'h3 ? _GEN_1148 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1251 = lvlReg == 2'h3 ? _GEN_1149 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1252 = lvlReg == 2'h3 ? _GEN_1150 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1253 = lvlReg == 2'h3 ? _GEN_1151 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1254 = lvlReg == 2'h3 ? _GEN_1152 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1255 = lvlReg == 2'h3 ? _GEN_1153 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1256 = lvlReg == 2'h3 ? _GEN_1154 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1257 = lvlReg == 2'h3 ? _GEN_1155 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1258 = lvlReg == 2'h3 ? _GEN_1156 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1259 = lvlReg == 2'h3 ? _GEN_1157 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1260 = lvlReg == 2'h3 ? _GEN_1158 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1261 = lvlReg == 2'h3 ? _GEN_1159 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1262 = lvlReg == 2'h3 ? _GEN_1160 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1263 = lvlReg == 2'h3 ? _GEN_1161 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1264 = lvlReg == 2'h3 ? _GEN_1162 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1265 = lvlReg == 2'h3 ? _GEN_1163 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1266 = lvlReg == 2'h3 ? _GEN_1164 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1267 = lvlReg == 2'h3 ? _GEN_1165 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1268 = lvlReg == 2'h3 ? _GEN_1166 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1269 = lvlReg == 2'h3 ? _GEN_1167 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1270 = lvlReg == 2'h3 ? _GEN_1168 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1271 = lvlReg == 2'h3 ? _GEN_1169 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1275 = lvlReg == 2'h3 ? _GEN_1173 : _GEN_195; // @[\\src\\main\\scala\\GameLogic.scala 478:34]
  wire  _GEN_1276 = lvlReg == 2'h3 ? _GEN_1174 : _GEN_196; // @[\\src\\main\\scala\\GameLogic.scala 478:34]
  wire  _GEN_1277 = lvlReg == 2'h3 ? _GEN_1175 : _GEN_197; // @[\\src\\main\\scala\\GameLogic.scala 478:34]
  wire  _GEN_1278 = lvlReg == 2'h3 ? _GEN_1176 : spriteVisibleRegs_64; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1279 = lvlReg == 2'h3 ? _GEN_1177 : spriteVisibleRegs_65; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1280 = lvlReg == 2'h3 ? _GEN_1178 : spriteVisibleRegs_66; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1281 = lvlReg == 2'h3 ? _GEN_1179 : spriteVisibleRegs_67; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1282 = lvlReg == 2'h3 ? _GEN_1180 : spriteVisibleRegs_68; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1283 = lvlReg == 2'h3 ? _GEN_1181 : spriteVisibleRegs_69; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1284 = lvlReg == 2'h3 ? _GEN_1182 : spriteVisibleRegs_70; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1285 = lvlReg == 2'h3 ? _GEN_1183 : spriteVisibleRegs_71; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1286 = lvlReg == 2'h3 ? _GEN_1184 : spriteVisibleRegs_72; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1287 = lvlReg == 2'h3 ? _GEN_1185 : spriteVisibleRegs_73; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1288 = lvlReg == 2'h3 ? _GEN_1186 : spriteVisibleRegs_74; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1289 = lvlReg == 2'h3 ? _GEN_1187 : spriteVisibleRegs_75; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1290 = lvlReg == 2'h3 ? _GEN_1188 : spriteVisibleRegs_76; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1291 = lvlReg == 2'h3 ? _GEN_1189 : spriteVisibleRegs_77; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1292 = lvlReg == 2'h3 ? _GEN_1190 : spriteVisibleRegs_78; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1293 = lvlReg == 2'h3 ? _GEN_1191 : spriteVisibleRegs_79; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1294 = lvlReg == 2'h3 ? _GEN_1192 : spriteVisibleRegs_80; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1295 = lvlReg == 2'h3 ? _GEN_1193 : spriteVisibleRegs_81; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1296 = lvlReg == 2'h3 ? _GEN_1194 : spriteVisibleRegs_82; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1297 = lvlReg == 2'h3 ? _GEN_1195 : spriteVisibleRegs_83; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1298 = lvlReg == 2'h3 ? _GEN_1196 : spriteVisibleRegs_84; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1299 = lvlReg == 2'h3 ? _GEN_1197 : spriteVisibleRegs_85; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1300 = lvlReg == 2'h3 ? _GEN_1198 : spriteVisibleRegs_86; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1301 = lvlReg == 2'h3 ? _GEN_1199 : spriteVisibleRegs_87; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1302 = lvlReg == 2'h3 ? _GEN_1200 : spriteVisibleRegs_88; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1303 = lvlReg == 2'h3 ? _GEN_1201 : spriteVisibleRegs_89; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1304 = lvlReg == 2'h3 ? _GEN_1202 : spriteVisibleRegs_90; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1305 = lvlReg == 2'h3 ? _GEN_1203 : spriteVisibleRegs_91; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1306 = lvlReg == 2'h3 ? _GEN_1204 : spriteVisibleRegs_92; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1307 = lvlReg == 2'h3 ? _GEN_1205 : spriteVisibleRegs_93; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1308 = lvlReg == 2'h3 ? _GEN_1206 : spriteVisibleRegs_94; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1309 = lvlReg == 2'h3 ? _GEN_1207 : spriteVisibleRegs_95; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1310 = lvlReg == 2'h3 ? _GEN_1208 : spriteVisibleRegs_96; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1311 = lvlReg == 2'h3 ? _GEN_1209 : spriteVisibleRegs_97; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1312 = lvlReg == 2'h3 ? _GEN_1210 : spriteVisibleRegs_98; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire  _GEN_1313 = lvlReg == 2'h3 ? _GEN_1211 : spriteVisibleRegs_99; // @[\\src\\main\\scala\\GameLogic.scala 125:34 478:34]
  wire [5:0] _GEN_1314 = lvlReg == 2'h3 ? _GEN_806 : nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 244:34 478:34]
  wire [7:0] _GEN_1315 = lvlReg == 2'h3 ? _GEN_1213 : spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 243:34 478:34]
  wire  _GEN_1319 = lvlReg == 2'h2 ? _GEN_912 : _GEN_1217; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1320 = lvlReg == 2'h2 ? _GEN_913 : _GEN_1218; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1321 = lvlReg == 2'h2 ? _GEN_914 : _GEN_1219; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1322 = lvlReg == 2'h2 ? _GEN_915 : _GEN_1220; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1323 = lvlReg == 2'h2 ? _GEN_916 : _GEN_1221; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1324 = lvlReg == 2'h2 ? _GEN_917 : _GEN_1222; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1325 = lvlReg == 2'h2 ? _GEN_918 : _GEN_1223; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1326 = lvlReg == 2'h2 ? _GEN_919 : _GEN_1224; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1327 = lvlReg == 2'h2 ? _GEN_920 : _GEN_1225; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1328 = lvlReg == 2'h2 ? _GEN_921 : _GEN_1226; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1329 = lvlReg == 2'h2 ? _GEN_922 : _GEN_1227; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1330 = lvlReg == 2'h2 ? _GEN_923 : _GEN_1228; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1331 = lvlReg == 2'h2 ? _GEN_924 : _GEN_1229; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1332 = lvlReg == 2'h2 ? _GEN_925 : _GEN_1230; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1333 = lvlReg == 2'h2 ? _GEN_926 : _GEN_1231; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1334 = lvlReg == 2'h2 ? _GEN_927 : _GEN_1232; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1335 = lvlReg == 2'h2 ? _GEN_928 : _GEN_1233; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1336 = lvlReg == 2'h2 ? _GEN_929 : _GEN_1234; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1337 = lvlReg == 2'h2 ? _GEN_930 : _GEN_1235; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1338 = lvlReg == 2'h2 ? _GEN_931 : _GEN_1236; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1339 = lvlReg == 2'h2 ? _GEN_932 : _GEN_1237; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1340 = lvlReg == 2'h2 ? _GEN_933 : _GEN_1238; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1341 = lvlReg == 2'h2 ? _GEN_934 : _GEN_1239; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1342 = lvlReg == 2'h2 ? _GEN_935 : _GEN_1240; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1343 = lvlReg == 2'h2 ? _GEN_936 : _GEN_1241; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1344 = lvlReg == 2'h2 ? _GEN_937 : _GEN_1242; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1345 = lvlReg == 2'h2 ? _GEN_938 : _GEN_1243; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1346 = lvlReg == 2'h2 ? _GEN_939 : _GEN_1244; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1347 = lvlReg == 2'h2 ? _GEN_940 : _GEN_1245; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1348 = lvlReg == 2'h2 ? _GEN_941 : _GEN_1246; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1349 = lvlReg == 2'h2 ? _GEN_942 : _GEN_1247; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1350 = lvlReg == 2'h2 ? _GEN_943 : _GEN_1248; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1351 = lvlReg == 2'h2 ? _GEN_944 : _GEN_1249; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1352 = lvlReg == 2'h2 ? _GEN_945 : _GEN_1250; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1353 = lvlReg == 2'h2 ? _GEN_946 : _GEN_1251; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1354 = lvlReg == 2'h2 ? _GEN_947 : _GEN_1252; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1355 = lvlReg == 2'h2 ? _GEN_948 : _GEN_1253; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1356 = lvlReg == 2'h2 ? _GEN_949 : _GEN_1254; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1357 = lvlReg == 2'h2 ? _GEN_950 : _GEN_1255; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1358 = lvlReg == 2'h2 ? _GEN_951 : _GEN_1256; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1359 = lvlReg == 2'h2 ? _GEN_952 : _GEN_1257; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1360 = lvlReg == 2'h2 ? _GEN_953 : _GEN_1258; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1361 = lvlReg == 2'h2 ? _GEN_954 : _GEN_1259; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1362 = lvlReg == 2'h2 ? _GEN_955 : _GEN_1260; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1363 = lvlReg == 2'h2 ? _GEN_956 : _GEN_1261; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1364 = lvlReg == 2'h2 ? _GEN_957 : _GEN_1262; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1365 = lvlReg == 2'h2 ? _GEN_958 : _GEN_1263; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1366 = lvlReg == 2'h2 ? _GEN_959 : _GEN_1264; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1367 = lvlReg == 2'h2 ? _GEN_960 : _GEN_1265; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1368 = lvlReg == 2'h2 ? _GEN_961 : _GEN_1266; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1369 = lvlReg == 2'h2 ? _GEN_962 : _GEN_1267; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1370 = lvlReg == 2'h2 ? _GEN_963 : _GEN_1268; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1371 = lvlReg == 2'h2 ? _GEN_964 : _GEN_1269; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1372 = lvlReg == 2'h2 ? _GEN_965 : _GEN_1270; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1373 = lvlReg == 2'h2 ? _GEN_966 : _GEN_1271; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1377 = lvlReg == 2'h2 ? _GEN_970 : _GEN_1275; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1378 = lvlReg == 2'h2 ? _GEN_971 : _GEN_1276; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1379 = lvlReg == 2'h2 ? _GEN_972 : _GEN_1277; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1380 = lvlReg == 2'h2 ? _GEN_973 : _GEN_1278; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1381 = lvlReg == 2'h2 ? _GEN_974 : _GEN_1279; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1382 = lvlReg == 2'h2 ? _GEN_975 : _GEN_1280; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1383 = lvlReg == 2'h2 ? _GEN_976 : _GEN_1281; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1384 = lvlReg == 2'h2 ? _GEN_977 : _GEN_1282; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1385 = lvlReg == 2'h2 ? _GEN_978 : _GEN_1283; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1386 = lvlReg == 2'h2 ? _GEN_979 : _GEN_1284; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1387 = lvlReg == 2'h2 ? _GEN_980 : _GEN_1285; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1388 = lvlReg == 2'h2 ? _GEN_981 : _GEN_1286; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1389 = lvlReg == 2'h2 ? _GEN_982 : _GEN_1287; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1390 = lvlReg == 2'h2 ? _GEN_983 : _GEN_1288; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1391 = lvlReg == 2'h2 ? _GEN_984 : _GEN_1289; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1392 = lvlReg == 2'h2 ? _GEN_985 : _GEN_1290; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1393 = lvlReg == 2'h2 ? _GEN_986 : _GEN_1291; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1394 = lvlReg == 2'h2 ? _GEN_987 : _GEN_1292; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1395 = lvlReg == 2'h2 ? _GEN_988 : _GEN_1293; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1396 = lvlReg == 2'h2 ? _GEN_989 : _GEN_1294; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1397 = lvlReg == 2'h2 ? _GEN_990 : _GEN_1295; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1398 = lvlReg == 2'h2 ? _GEN_991 : _GEN_1296; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1399 = lvlReg == 2'h2 ? _GEN_992 : _GEN_1297; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1400 = lvlReg == 2'h2 ? _GEN_993 : _GEN_1298; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1401 = lvlReg == 2'h2 ? _GEN_994 : _GEN_1299; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1402 = lvlReg == 2'h2 ? _GEN_995 : _GEN_1300; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1403 = lvlReg == 2'h2 ? _GEN_996 : _GEN_1301; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1404 = lvlReg == 2'h2 ? _GEN_997 : _GEN_1302; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1405 = lvlReg == 2'h2 ? _GEN_998 : _GEN_1303; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1406 = lvlReg == 2'h2 ? _GEN_999 : _GEN_1304; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1407 = lvlReg == 2'h2 ? _GEN_1000 : _GEN_1305; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1408 = lvlReg == 2'h2 ? _GEN_1001 : _GEN_1306; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1409 = lvlReg == 2'h2 ? _GEN_1002 : _GEN_1307; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1410 = lvlReg == 2'h2 ? _GEN_1003 : _GEN_1308; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1411 = lvlReg == 2'h2 ? _GEN_1004 : _GEN_1309; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1412 = lvlReg == 2'h2 ? _GEN_1005 : _GEN_1310; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1413 = lvlReg == 2'h2 ? _GEN_1006 : _GEN_1311; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1414 = lvlReg == 2'h2 ? _GEN_1007 : _GEN_1312; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1415 = lvlReg == 2'h2 ? _GEN_1008 : _GEN_1313; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire [5:0] _GEN_1416 = lvlReg == 2'h2 ? _GEN_806 : _GEN_1314; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire [7:0] _GEN_1417 = lvlReg == 2'h2 ? _GEN_1010 : _GEN_1315; // @[\\src\\main\\scala\\GameLogic.scala 469:34]
  wire  _GEN_1431 = lvlReg == 2'h1 ? _GEN_719 : _GEN_1329; // @[\\src\\main\\scala\\GameLogic.scala 460:28]
  wire  _GEN_1432 = lvlReg == 2'h1 ? _GEN_720 : _GEN_1330; // @[\\src\\main\\scala\\GameLogic.scala 460:28]
  wire  _T_90 = ~isBlinking; // @[\\src\\main\\scala\\GameLogic.scala 492:12]
  wire [6:0] _obstacleWidth_T_1 = 5'h1a * 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 497:81]
  wire [5:0] _obstacleHeight_T_1 = 4'hf * 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 498:83]
  wire [6:0] _T_93 = spriteScaleTypeRegs_0 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2715 = {{4{_T_93[6]}},_T_93}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_96 = $signed(spriteXRegs_16) + $signed(_GEN_2715); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_97 = $signed(spriteXRegs_14) < $signed(_T_96); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_98 = spriteVisibleRegs_16 & $signed(spriteXRegs_16) <= 11'sh280 & _T_97; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [10:0] _T_101 = $signed(spriteXRegs_14) + 11'sh8; // @[\\src\\main\\scala\\GameLogic.scala 502:110]
  wire [5:0] _T_104 = spriteScaleTypeRegs_0 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2716 = {{4{_T_104[5]}},_T_104}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_107 = $signed(spriteYRegs_16) + $signed(_GEN_2716); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_108 = $signed(spriteYRegs_14) < $signed(_T_107); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_109 = _T_98 & $signed(spriteXRegs_16) < $signed(_T_101) & _T_108; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire [9:0] _T_112 = $signed(spriteYRegs_14) + 10'shb; // @[\\src\\main\\scala\\GameLogic.scala 503:111]
  wire  _T_114 = _T_109 & $signed(spriteYRegs_16) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire  _GEN_1520 = _T_114 | collisionDetected; // @[\\src\\main\\scala\\GameLogic.scala 504:13 505:31 250:34]
  wire [6:0] _T_117 = spriteScaleTypeRegs_1 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2717 = {{4{_T_117[6]}},_T_117}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_120 = $signed(spriteXRegs_17) + $signed(_GEN_2717); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_121 = $signed(spriteXRegs_14) < $signed(_T_120); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_122 = spriteVisibleRegs_17 & $signed(spriteXRegs_17) <= 11'sh280 & _T_121; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [5:0] _T_128 = spriteScaleTypeRegs_1 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2718 = {{4{_T_128[5]}},_T_128}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_131 = $signed(spriteYRegs_17) + $signed(_GEN_2718); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_132 = $signed(spriteYRegs_14) < $signed(_T_131); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_133 = _T_122 & $signed(spriteXRegs_17) < $signed(_T_101) & _T_132; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire  _T_138 = _T_133 & $signed(spriteYRegs_17) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire [6:0] _T_141 = spriteScaleTypeRegs_2 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2719 = {{4{_T_141[6]}},_T_141}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_144 = $signed(spriteXRegs_18) + $signed(_GEN_2719); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_145 = $signed(spriteXRegs_14) < $signed(_T_144); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_146 = spriteVisibleRegs_18 & $signed(spriteXRegs_18) <= 11'sh280 & _T_145; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [5:0] _T_152 = spriteScaleTypeRegs_2 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2720 = {{4{_T_152[5]}},_T_152}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_155 = $signed(spriteYRegs_18) + $signed(_GEN_2720); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_156 = $signed(spriteYRegs_14) < $signed(_T_155); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_157 = _T_146 & $signed(spriteXRegs_18) < $signed(_T_101) & _T_156; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire  _T_162 = _T_157 & $signed(spriteYRegs_18) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire [6:0] _T_165 = spriteScaleTypeRegs_3 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2721 = {{4{_T_165[6]}},_T_165}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_168 = $signed(spriteXRegs_19) + $signed(_GEN_2721); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_169 = $signed(spriteXRegs_14) < $signed(_T_168); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_170 = spriteVisibleRegs_19 & $signed(spriteXRegs_19) <= 11'sh280 & _T_169; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [5:0] _T_176 = spriteScaleTypeRegs_3 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2722 = {{4{_T_176[5]}},_T_176}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_179 = $signed(spriteYRegs_19) + $signed(_GEN_2722); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_180 = $signed(spriteYRegs_14) < $signed(_T_179); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_181 = _T_170 & $signed(spriteXRegs_19) < $signed(_T_101) & _T_180; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire  _T_186 = _T_181 & $signed(spriteYRegs_19) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire [6:0] _T_189 = spriteScaleTypeRegs_4 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2723 = {{4{_T_189[6]}},_T_189}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_192 = $signed(spriteXRegs_20) + $signed(_GEN_2723); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_193 = $signed(spriteXRegs_14) < $signed(_T_192); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_194 = spriteVisibleRegs_20 & $signed(spriteXRegs_20) <= 11'sh280 & _T_193; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [5:0] _T_200 = spriteScaleTypeRegs_4 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2724 = {{4{_T_200[5]}},_T_200}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_203 = $signed(spriteYRegs_20) + $signed(_GEN_2724); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_204 = $signed(spriteYRegs_14) < $signed(_T_203); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_205 = _T_194 & $signed(spriteXRegs_20) < $signed(_T_101) & _T_204; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire  _T_210 = _T_205 & $signed(spriteYRegs_20) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire [6:0] _T_213 = spriteScaleTypeRegs_5 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2725 = {{4{_T_213[6]}},_T_213}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_216 = $signed(spriteXRegs_21) + $signed(_GEN_2725); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_217 = $signed(spriteXRegs_14) < $signed(_T_216); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_218 = spriteVisibleRegs_21 & $signed(spriteXRegs_21) <= 11'sh280 & _T_217; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [5:0] _T_224 = spriteScaleTypeRegs_5 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2726 = {{4{_T_224[5]}},_T_224}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_227 = $signed(spriteYRegs_21) + $signed(_GEN_2726); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_228 = $signed(spriteYRegs_14) < $signed(_T_227); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_229 = _T_218 & $signed(spriteXRegs_21) < $signed(_T_101) & _T_228; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire  _T_234 = _T_229 & $signed(spriteYRegs_21) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire [6:0] _T_237 = spriteScaleTypeRegs_6 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2727 = {{4{_T_237[6]}},_T_237}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_240 = $signed(spriteXRegs_22) + $signed(_GEN_2727); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_241 = $signed(spriteXRegs_14) < $signed(_T_240); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_242 = spriteVisibleRegs_22 & $signed(spriteXRegs_22) <= 11'sh280 & _T_241; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [5:0] _T_248 = spriteScaleTypeRegs_6 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2728 = {{4{_T_248[5]}},_T_248}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_251 = $signed(spriteYRegs_22) + $signed(_GEN_2728); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_252 = $signed(spriteYRegs_14) < $signed(_T_251); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_253 = _T_242 & $signed(spriteXRegs_22) < $signed(_T_101) & _T_252; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire  _T_258 = _T_253 & $signed(spriteYRegs_22) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire [6:0] _T_261 = spriteScaleTypeRegs_7 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2729 = {{4{_T_261[6]}},_T_261}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_264 = $signed(spriteXRegs_23) + $signed(_GEN_2729); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_265 = $signed(spriteXRegs_14) < $signed(_T_264); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_266 = spriteVisibleRegs_23 & $signed(spriteXRegs_23) <= 11'sh280 & _T_265; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [5:0] _T_272 = spriteScaleTypeRegs_7 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2730 = {{4{_T_272[5]}},_T_272}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_275 = $signed(spriteYRegs_23) + $signed(_GEN_2730); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_276 = $signed(spriteYRegs_14) < $signed(_T_275); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_277 = _T_266 & $signed(spriteXRegs_23) < $signed(_T_101) & _T_276; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire  _T_282 = _T_277 & $signed(spriteYRegs_23) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire [6:0] _T_285 = spriteScaleTypeRegs_8 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2731 = {{4{_T_285[6]}},_T_285}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_288 = $signed(spriteXRegs_24) + $signed(_GEN_2731); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_289 = $signed(spriteXRegs_14) < $signed(_T_288); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_290 = spriteVisibleRegs_24 & $signed(spriteXRegs_24) <= 11'sh280 & _T_289; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [5:0] _T_296 = spriteScaleTypeRegs_8 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2732 = {{4{_T_296[5]}},_T_296}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_299 = $signed(spriteYRegs_24) + $signed(_GEN_2732); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_300 = $signed(spriteYRegs_14) < $signed(_T_299); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_301 = _T_290 & $signed(spriteXRegs_24) < $signed(_T_101) & _T_300; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire  _T_306 = _T_301 & $signed(spriteYRegs_24) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire [6:0] _T_309 = spriteScaleTypeRegs_9 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 502:65]
  wire [10:0] _GEN_2733 = {{4{_T_309[6]}},_T_309}; // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire [10:0] _T_312 = $signed(spriteXRegs_25) + $signed(_GEN_2733); // @[\\src\\main\\scala\\GameLogic.scala 502:49]
  wire  _T_313 = $signed(spriteXRegs_14) < $signed(_T_312); // @[\\src\\main\\scala\\GameLogic.scala 502:32]
  wire  _T_314 = spriteVisibleRegs_25 & $signed(spriteXRegs_25) <= 11'sh280 & _T_313; // @[\\src\\main\\scala\\GameLogic.scala 501:63]
  wire [5:0] _T_320 = spriteScaleTypeRegs_9 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 503:66]
  wire [9:0] _GEN_2734 = {{4{_T_320[5]}},_T_320}; // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire [9:0] _T_323 = $signed(spriteYRegs_25) + $signed(_GEN_2734); // @[\\src\\main\\scala\\GameLogic.scala 503:49]
  wire  _T_324 = $signed(spriteYRegs_14) < $signed(_T_323); // @[\\src\\main\\scala\\GameLogic.scala 503:32]
  wire  _T_325 = _T_314 & $signed(spriteXRegs_25) < $signed(_T_101) & _T_324; // @[\\src\\main\\scala\\GameLogic.scala 502:117]
  wire  _T_330 = _T_325 & $signed(spriteYRegs_25) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 503:74]
  wire  _GEN_1529 = _T_330 | (_T_306 | (_T_282 | (_T_258 | (_T_234 | (_T_210 | (_T_186 | (_T_162 | (_T_138 | _GEN_1520))
    )))))); // @[\\src\\main\\scala\\GameLogic.scala 504:13 505:31]
  wire  _GEN_1530 = ~isBlinking ? _GEN_1529 : collisionDetected; // @[\\src\\main\\scala\\GameLogic.scala 492:25 250:34]
  wire [6:0] _obstacleWidth_T_21 = 5'h1d * 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 515:81]
  wire [6:0] _T_332 = spriteScaleTypeRegs_0 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2735 = {{4{_T_332[6]}},_T_332}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_335 = $signed(spriteXRegs_26) + $signed(_GEN_2735); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_336 = $signed(spriteXRegs_14) < $signed(_T_335); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_337 = spriteVisibleRegs_26 & _T_336; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_346 = $signed(spriteYRegs_26) + $signed(_GEN_2716); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_347 = $signed(spriteYRegs_14) < $signed(_T_346); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_348 = _T_337 & $signed(spriteXRegs_26) < $signed(_T_101) & _T_347; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_353 = _T_348 & $signed(spriteYRegs_26) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire [6:0] _T_354 = spriteScaleTypeRegs_1 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2737 = {{4{_T_354[6]}},_T_354}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_357 = $signed(spriteXRegs_27) + $signed(_GEN_2737); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_358 = $signed(spriteXRegs_14) < $signed(_T_357); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_359 = spriteVisibleRegs_27 & _T_358; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_368 = $signed(spriteYRegs_27) + $signed(_GEN_2718); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_369 = $signed(spriteYRegs_14) < $signed(_T_368); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_370 = _T_359 & $signed(spriteXRegs_27) < $signed(_T_101) & _T_369; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_375 = _T_370 & $signed(spriteYRegs_27) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire [6:0] _T_376 = spriteScaleTypeRegs_2 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2739 = {{4{_T_376[6]}},_T_376}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_379 = $signed(spriteXRegs_28) + $signed(_GEN_2739); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_380 = $signed(spriteXRegs_14) < $signed(_T_379); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_381 = spriteVisibleRegs_28 & _T_380; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_390 = $signed(spriteYRegs_28) + $signed(_GEN_2720); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_391 = $signed(spriteYRegs_14) < $signed(_T_390); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_392 = _T_381 & $signed(spriteXRegs_28) < $signed(_T_101) & _T_391; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_397 = _T_392 & $signed(spriteYRegs_28) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire [6:0] _T_398 = spriteScaleTypeRegs_3 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2741 = {{4{_T_398[6]}},_T_398}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_401 = $signed(spriteXRegs_29) + $signed(_GEN_2741); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_402 = $signed(spriteXRegs_14) < $signed(_T_401); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_403 = spriteVisibleRegs_29 & _T_402; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_412 = $signed(spriteYRegs_29) + $signed(_GEN_2722); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_413 = $signed(spriteYRegs_14) < $signed(_T_412); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_414 = _T_403 & $signed(spriteXRegs_29) < $signed(_T_101) & _T_413; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_419 = _T_414 & $signed(spriteYRegs_29) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire [6:0] _T_420 = spriteScaleTypeRegs_4 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2743 = {{4{_T_420[6]}},_T_420}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_423 = $signed(spriteXRegs_30) + $signed(_GEN_2743); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_424 = $signed(spriteXRegs_14) < $signed(_T_423); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_425 = spriteVisibleRegs_30 & _T_424; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_434 = $signed(spriteYRegs_30) + $signed(_GEN_2724); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_435 = $signed(spriteYRegs_14) < $signed(_T_434); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_436 = _T_425 & $signed(spriteXRegs_30) < $signed(_T_101) & _T_435; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_441 = _T_436 & $signed(spriteYRegs_30) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire [6:0] _T_442 = spriteScaleTypeRegs_5 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2745 = {{4{_T_442[6]}},_T_442}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_445 = $signed(spriteXRegs_31) + $signed(_GEN_2745); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_446 = $signed(spriteXRegs_14) < $signed(_T_445); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_447 = spriteVisibleRegs_31 & _T_446; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_456 = $signed(spriteYRegs_31) + $signed(_GEN_2726); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_457 = $signed(spriteYRegs_14) < $signed(_T_456); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_458 = _T_447 & $signed(spriteXRegs_31) < $signed(_T_101) & _T_457; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_463 = _T_458 & $signed(spriteYRegs_31) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire [6:0] _T_464 = spriteScaleTypeRegs_6 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2747 = {{4{_T_464[6]}},_T_464}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_467 = $signed(spriteXRegs_32) + $signed(_GEN_2747); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_468 = $signed(spriteXRegs_14) < $signed(_T_467); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_469 = spriteVisibleRegs_32 & _T_468; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_478 = $signed(spriteYRegs_32) + $signed(_GEN_2728); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_479 = $signed(spriteYRegs_14) < $signed(_T_478); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_480 = _T_469 & $signed(spriteXRegs_32) < $signed(_T_101) & _T_479; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_485 = _T_480 & $signed(spriteYRegs_32) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire [6:0] _T_486 = spriteScaleTypeRegs_7 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2749 = {{4{_T_486[6]}},_T_486}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_489 = $signed(spriteXRegs_33) + $signed(_GEN_2749); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_490 = $signed(spriteXRegs_14) < $signed(_T_489); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_491 = spriteVisibleRegs_33 & _T_490; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_500 = $signed(spriteYRegs_33) + $signed(_GEN_2730); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_501 = $signed(spriteYRegs_14) < $signed(_T_500); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_502 = _T_491 & $signed(spriteXRegs_33) < $signed(_T_101) & _T_501; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_507 = _T_502 & $signed(spriteYRegs_33) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire [6:0] _T_508 = spriteScaleTypeRegs_8 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2751 = {{4{_T_508[6]}},_T_508}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_511 = $signed(spriteXRegs_34) + $signed(_GEN_2751); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_512 = $signed(spriteXRegs_14) < $signed(_T_511); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_513 = spriteVisibleRegs_34 & _T_512; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_522 = $signed(spriteYRegs_34) + $signed(_GEN_2732); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_523 = $signed(spriteYRegs_14) < $signed(_T_522); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_524 = _T_513 & $signed(spriteXRegs_34) < $signed(_T_101) & _T_523; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_529 = _T_524 & $signed(spriteYRegs_34) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire [6:0] _T_530 = spriteScaleTypeRegs_9 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 520:65]
  wire [10:0] _GEN_2753 = {{4{_T_530[6]}},_T_530}; // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire [10:0] _T_533 = $signed(spriteXRegs_35) + $signed(_GEN_2753); // @[\\src\\main\\scala\\GameLogic.scala 520:49]
  wire  _T_534 = $signed(spriteXRegs_14) < $signed(_T_533); // @[\\src\\main\\scala\\GameLogic.scala 520:32]
  wire  _T_535 = spriteVisibleRegs_35 & _T_534; // @[\\src\\main\\scala\\GameLogic.scala 519:34]
  wire [9:0] _T_544 = $signed(spriteYRegs_35) + $signed(_GEN_2734); // @[\\src\\main\\scala\\GameLogic.scala 521:49]
  wire  _T_545 = $signed(spriteYRegs_14) < $signed(_T_544); // @[\\src\\main\\scala\\GameLogic.scala 521:32]
  wire  _T_546 = _T_535 & $signed(spriteXRegs_35) < $signed(_T_101) & _T_545; // @[\\src\\main\\scala\\GameLogic.scala 520:117]
  wire  _T_551 = _T_546 & $signed(spriteYRegs_35) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 521:74]
  wire  _GEN_1540 = _T_551 | (_T_529 | (_T_507 | (_T_485 | (_T_463 | (_T_441 | (_T_419 | (_T_397 | (_T_375 | (_T_353 |
    _GEN_1530))))))))); // @[\\src\\main\\scala\\GameLogic.scala 522:13 523:31]
  wire  _GEN_1541 = _T_90 ? _GEN_1540 : _GEN_1530; // @[\\src\\main\\scala\\GameLogic.scala 510:25]
  wire [7:0] _obstacleWidth_T_41 = 6'h20 * 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 533:81]
  wire [7:0] _T_553 = spriteScaleTypeRegs_0 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2755 = {{3{_T_553[7]}},_T_553}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_556 = $signed(spriteXRegs_36) + $signed(_GEN_2755); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_557 = $signed(spriteXRegs_14) < $signed(_T_556); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_558 = spriteVisibleRegs_36 & _T_557; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_567 = $signed(spriteYRegs_36) + $signed(_GEN_2716); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_568 = $signed(spriteYRegs_14) < $signed(_T_567); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_569 = _T_558 & $signed(spriteXRegs_36) < $signed(_T_101) & _T_568; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_574 = _T_569 & $signed(spriteYRegs_36) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire [7:0] _T_575 = spriteScaleTypeRegs_1 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2757 = {{3{_T_575[7]}},_T_575}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_578 = $signed(spriteXRegs_37) + $signed(_GEN_2757); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_579 = $signed(spriteXRegs_14) < $signed(_T_578); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_580 = spriteVisibleRegs_37 & _T_579; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_589 = $signed(spriteYRegs_37) + $signed(_GEN_2718); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_590 = $signed(spriteYRegs_14) < $signed(_T_589); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_591 = _T_580 & $signed(spriteXRegs_37) < $signed(_T_101) & _T_590; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_596 = _T_591 & $signed(spriteYRegs_37) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire [7:0] _T_597 = spriteScaleTypeRegs_2 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2759 = {{3{_T_597[7]}},_T_597}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_600 = $signed(spriteXRegs_38) + $signed(_GEN_2759); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_601 = $signed(spriteXRegs_14) < $signed(_T_600); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_602 = spriteVisibleRegs_38 & _T_601; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_611 = $signed(spriteYRegs_38) + $signed(_GEN_2720); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_612 = $signed(spriteYRegs_14) < $signed(_T_611); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_613 = _T_602 & $signed(spriteXRegs_38) < $signed(_T_101) & _T_612; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_618 = _T_613 & $signed(spriteYRegs_38) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire [7:0] _T_619 = spriteScaleTypeRegs_3 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2761 = {{3{_T_619[7]}},_T_619}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_622 = $signed(spriteXRegs_39) + $signed(_GEN_2761); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_623 = $signed(spriteXRegs_14) < $signed(_T_622); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_624 = spriteVisibleRegs_39 & _T_623; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_633 = $signed(spriteYRegs_39) + $signed(_GEN_2722); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_634 = $signed(spriteYRegs_14) < $signed(_T_633); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_635 = _T_624 & $signed(spriteXRegs_39) < $signed(_T_101) & _T_634; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_640 = _T_635 & $signed(spriteYRegs_39) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire [7:0] _T_641 = spriteScaleTypeRegs_4 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2763 = {{3{_T_641[7]}},_T_641}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_644 = $signed(spriteXRegs_40) + $signed(_GEN_2763); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_645 = $signed(spriteXRegs_14) < $signed(_T_644); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_646 = spriteVisibleRegs_40 & _T_645; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_655 = $signed(spriteYRegs_40) + $signed(_GEN_2724); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_656 = $signed(spriteYRegs_14) < $signed(_T_655); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_657 = _T_646 & $signed(spriteXRegs_40) < $signed(_T_101) & _T_656; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_662 = _T_657 & $signed(spriteYRegs_40) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire [7:0] _T_663 = spriteScaleTypeRegs_5 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2765 = {{3{_T_663[7]}},_T_663}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_666 = $signed(spriteXRegs_41) + $signed(_GEN_2765); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_667 = $signed(spriteXRegs_14) < $signed(_T_666); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_668 = spriteVisibleRegs_41 & _T_667; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_677 = $signed(spriteYRegs_41) + $signed(_GEN_2726); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_678 = $signed(spriteYRegs_14) < $signed(_T_677); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_679 = _T_668 & $signed(spriteXRegs_41) < $signed(_T_101) & _T_678; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_684 = _T_679 & $signed(spriteYRegs_41) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire [7:0] _T_685 = spriteScaleTypeRegs_6 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2767 = {{3{_T_685[7]}},_T_685}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_688 = $signed(spriteXRegs_42) + $signed(_GEN_2767); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_689 = $signed(spriteXRegs_14) < $signed(_T_688); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_690 = spriteVisibleRegs_42 & _T_689; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_699 = $signed(spriteYRegs_42) + $signed(_GEN_2728); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_700 = $signed(spriteYRegs_14) < $signed(_T_699); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_701 = _T_690 & $signed(spriteXRegs_42) < $signed(_T_101) & _T_700; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_706 = _T_701 & $signed(spriteYRegs_42) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire [7:0] _T_707 = spriteScaleTypeRegs_7 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2769 = {{3{_T_707[7]}},_T_707}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_710 = $signed(spriteXRegs_43) + $signed(_GEN_2769); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_711 = $signed(spriteXRegs_14) < $signed(_T_710); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_712 = spriteVisibleRegs_43 & _T_711; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_721 = $signed(spriteYRegs_43) + $signed(_GEN_2730); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_722 = $signed(spriteYRegs_14) < $signed(_T_721); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_723 = _T_712 & $signed(spriteXRegs_43) < $signed(_T_101) & _T_722; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_728 = _T_723 & $signed(spriteYRegs_43) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire [7:0] _T_729 = spriteScaleTypeRegs_8 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2771 = {{3{_T_729[7]}},_T_729}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_732 = $signed(spriteXRegs_44) + $signed(_GEN_2771); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_733 = $signed(spriteXRegs_14) < $signed(_T_732); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_734 = spriteVisibleRegs_44 & _T_733; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_743 = $signed(spriteYRegs_44) + $signed(_GEN_2732); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_744 = $signed(spriteYRegs_14) < $signed(_T_743); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_745 = _T_734 & $signed(spriteXRegs_44) < $signed(_T_101) & _T_744; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_750 = _T_745 & $signed(spriteYRegs_44) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire [7:0] _T_751 = spriteScaleTypeRegs_9 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 537:65]
  wire [10:0] _GEN_2773 = {{3{_T_751[7]}},_T_751}; // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire [10:0] _T_754 = $signed(spriteXRegs_45) + $signed(_GEN_2773); // @[\\src\\main\\scala\\GameLogic.scala 537:49]
  wire  _T_755 = $signed(spriteXRegs_14) < $signed(_T_754); // @[\\src\\main\\scala\\GameLogic.scala 537:32]
  wire  _T_756 = spriteVisibleRegs_45 & _T_755; // @[\\src\\main\\scala\\GameLogic.scala 536:34]
  wire [9:0] _T_765 = $signed(spriteYRegs_45) + $signed(_GEN_2734); // @[\\src\\main\\scala\\GameLogic.scala 538:49]
  wire  _T_766 = $signed(spriteYRegs_14) < $signed(_T_765); // @[\\src\\main\\scala\\GameLogic.scala 538:32]
  wire  _T_767 = _T_756 & $signed(spriteXRegs_45) < $signed(_T_101) & _T_766; // @[\\src\\main\\scala\\GameLogic.scala 537:117]
  wire  _T_772 = _T_767 & $signed(spriteYRegs_45) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 538:74]
  wire  _GEN_1551 = _T_772 | (_T_750 | (_T_728 | (_T_706 | (_T_684 | (_T_662 | (_T_640 | (_T_618 | (_T_596 | (_T_574 |
    _GEN_1541))))))))); // @[\\src\\main\\scala\\GameLogic.scala 539:13 540:31]
  wire  _GEN_1552 = _T_90 ? _GEN_1551 : _GEN_1541; // @[\\src\\main\\scala\\GameLogic.scala 528:25]
  wire [10:0] _T_775 = $signed(spriteXRegs_13) + 11'sh16; // @[\\src\\main\\scala\\GameLogic.scala 548:46]
  wire  _T_776 = $signed(spriteXRegs_14) < $signed(_T_775); // @[\\src\\main\\scala\\GameLogic.scala 548:28]
  wire  _T_777 = spriteVisibleRegs_13 & _T_776; // @[\\src\\main\\scala\\GameLogic.scala 547:31]
  wire [9:0] _T_785 = $signed(spriteYRegs_13) + 10'sh16; // @[\\src\\main\\scala\\GameLogic.scala 549:46]
  wire  _T_786 = $signed(spriteYRegs_14) < $signed(_T_785); // @[\\src\\main\\scala\\GameLogic.scala 549:28]
  wire  _T_787 = _T_777 & $signed(spriteXRegs_13) < $signed(_T_101) & _T_786; // @[\\src\\main\\scala\\GameLogic.scala 548:99]
  wire  _T_792 = _T_787 & $signed(spriteYRegs_13) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 549:54]
  wire [2:0] _livesReg_T_1 = livesReg + 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 553:32]
  wire [2:0] _GEN_1553 = livesReg < 3'h3 ? _livesReg_T_1 : livesReg; // @[\\src\\main\\scala\\GameLogic.scala 552:30 553:20 231:25]
  wire [2:0] _GEN_1555 = _T_792 ? _GEN_1553 : livesReg; // @[\\src\\main\\scala\\GameLogic.scala 231:25 550:9]
  wire  _GEN_1556 = collisionDetected & _T_90 | isBlinking; // @[\\src\\main\\scala\\GameLogic.scala 558:46 559:20 253:27]
  wire [7:0] _GEN_1557 = collisionDetected & _T_90 ? 8'h0 : blinkCounter; // @[\\src\\main\\scala\\GameLogic.scala 558:46 560:22 251:29]
  wire [1:0] _GEN_1558 = collisionDetected & _T_90 ? 2'h0 : blinkTimes; // @[\\src\\main\\scala\\GameLogic.scala 558:46 561:20 252:27]
  wire  _GEN_1559 = blinkCounter < 8'h14 | _GEN_1432; // @[\\src\\main\\scala\\GameLogic.scala 569:41 570:33]
  wire  _GEN_1560 = blinkCounter < 8'ha ? 1'h0 : _GEN_1559; // @[\\src\\main\\scala\\GameLogic.scala 567:35 568:33]
  wire [7:0] _blinkCounter_T_1 = blinkCounter + 8'h1; // @[\\src\\main\\scala\\GameLogic.scala 572:38]
  wire [1:0] _blinkTimes_T_1 = blinkTimes + 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 575:36]
  wire [7:0] _GEN_1561 = blinkCounter == 8'h14 ? 8'h0 : _blinkCounter_T_1; // @[\\src\\main\\scala\\GameLogic.scala 572:22 573:37 574:24]
  wire [1:0] _GEN_1562 = blinkCounter == 8'h14 ? _blinkTimes_T_1 : _GEN_1558; // @[\\src\\main\\scala\\GameLogic.scala 573:37 575:22]
  wire [2:0] _livesReg_T_3 = livesReg - 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 584:34]
  wire [2:0] _GEN_1563 = livesReg <= 3'h1 ? 3'h0 : _livesReg_T_3; // @[\\src\\main\\scala\\GameLogic.scala 580:33 581:22 584:22]
  wire [2:0] _GEN_1564 = livesReg <= 3'h1 ? 3'h6 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 580:33 582:22 113:25]
  wire  _GEN_1565 = blinkTimes == 2'h3 ? 1'h0 : _GEN_1556; // @[\\src\\main\\scala\\GameLogic.scala 577:34 578:22]
  wire  _GEN_1566 = blinkTimes == 2'h3 | _GEN_1560; // @[\\src\\main\\scala\\GameLogic.scala 577:34 579:33]
  wire [2:0] _GEN_1567 = blinkTimes == 2'h3 ? _GEN_1563 : _GEN_1555; // @[\\src\\main\\scala\\GameLogic.scala 577:34]
  wire [2:0] _GEN_1568 = blinkTimes == 2'h3 ? _GEN_1564 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 113:25 577:34]
  wire  _GEN_1569 = blinkTimes == 2'h3 ? 1'h0 : _GEN_1552; // @[\\src\\main\\scala\\GameLogic.scala 577:34 586:29]
  wire [2:0] _GEN_1575 = isBlinking ? _GEN_1568 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 565:24 113:25]
  reg [10:0] spriteXRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 605:35]
  reg [9:0] spriteYRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 606:35]
  reg [10:0] spriteXRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 607:35]
  reg [9:0] spriteYRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 608:35]
  reg [10:0] spriteXRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 609:35]
  reg [9:0] spriteYRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 610:35]
  wire [9:0] _starCnt_T_1 = starCnt + 10'h1; // @[\\src\\main\\scala\\GameLogic.scala 617:28]
  wire [10:0] _spriteXRegs_58_T_5 = $signed(spriteXRegs_58) + 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 625:44]
  wire [10:0] _spriteXRegs_59_T_5 = $signed(spriteXRegs_59) + 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 626:44]
  wire [10:0] _spriteXRegs_60_T_5 = $signed(spriteXRegs_60) + 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 627:44]
  wire [9:0] _spriteYRegs_58_T_5 = $signed(spriteYRegs_58) + 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 628:44]
  wire [9:0] _spriteYRegs_59_T_5 = $signed(spriteYRegs_59) + 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 629:44]
  wire [9:0] _spriteYRegs_60_T_5 = $signed(spriteYRegs_60) + 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 630:44]
  reg [10:0] spriteXRegs_58_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 633:35]
  reg [9:0] spriteYRegs_58_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 634:35]
  reg [10:0] spriteXRegs_59_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 635:35]
  reg [9:0] spriteYRegs_59_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 636:35]
  reg [10:0] spriteXRegs_60_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 637:35]
  reg [9:0] spriteYRegs_60_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 638:35]
  reg [10:0] spriteXRegs_58_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 661:35]
  reg [9:0] spriteYRegs_58_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 662:35]
  reg [10:0] spriteXRegs_59_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 663:35]
  reg [9:0] spriteYRegs_59_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 664:35]
  reg [10:0] spriteXRegs_60_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 665:35]
  reg [9:0] spriteYRegs_60_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 666:35]
  wire [9:0] _GEN_1578 = starCnt == 10'h168 ? 10'h0 : _starCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 688:37 689:17 691:17]
  wire  _GEN_1579 = starCnt == 10'h12c ? 1'h0 : sprite58ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 674:37 675:35 176:42]
  wire  _GEN_1580 = starCnt == 10'h12c ? 1'h0 : sprite59ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 674:37 676:35 178:42]
  wire  _GEN_1581 = starCnt == 10'h12c ? 1'h0 : sprite60ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 674:37 677:35 180:42]
  wire  _GEN_1582 = starCnt == 10'h12c ? 1'h0 : sprite58ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 674:37 678:33 177:40]
  wire  _GEN_1583 = starCnt == 10'h12c ? 1'h0 : sprite59ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 674:37 679:33 179:40]
  wire  _GEN_1584 = starCnt == 10'h12c ? 1'h0 : sprite60ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 674:37 680:33 181:40]
  wire [10:0] _GEN_1585 = starCnt == 10'h12c ? $signed(_spriteXRegs_58_T_5) : $signed(_GEN_102); // @[\\src\\main\\scala\\GameLogic.scala 674:37 681:25]
  wire [10:0] _GEN_1586 = starCnt == 10'h12c ? $signed(_spriteXRegs_59_T_5) : $signed(_GEN_104); // @[\\src\\main\\scala\\GameLogic.scala 674:37 682:25]
  wire [10:0] _GEN_1587 = starCnt == 10'h12c ? $signed(_spriteXRegs_60_T_5) : $signed(_GEN_106); // @[\\src\\main\\scala\\GameLogic.scala 674:37 683:25]
  wire [9:0] _GEN_1588 = starCnt == 10'h12c ? $signed(_spriteYRegs_58_T_5) : $signed(_GEN_103); // @[\\src\\main\\scala\\GameLogic.scala 674:37 684:25]
  wire [9:0] _GEN_1589 = starCnt == 10'h12c ? $signed(_spriteYRegs_59_T_5) : $signed(_GEN_105); // @[\\src\\main\\scala\\GameLogic.scala 674:37 685:25]
  wire [9:0] _GEN_1590 = starCnt == 10'h12c ? $signed(_spriteYRegs_60_T_5) : $signed(_GEN_107); // @[\\src\\main\\scala\\GameLogic.scala 674:37 686:25]
  wire [9:0] _GEN_1591 = starCnt == 10'h12c ? _starCnt_T_1 : _GEN_1578; // @[\\src\\main\\scala\\GameLogic.scala 674:37 687:17]
  wire [10:0] _GEN_1592 = starCnt == 10'hf0 ? $signed(spriteXRegs_58_REG_2) : $signed(_GEN_1585); // @[\\src\\main\\scala\\GameLogic.scala 660:37 661:25]
  wire [9:0] _GEN_1593 = starCnt == 10'hf0 ? $signed(spriteYRegs_58_REG_2) : $signed(_GEN_1588); // @[\\src\\main\\scala\\GameLogic.scala 660:37 662:25]
  wire [10:0] _GEN_1594 = starCnt == 10'hf0 ? $signed(spriteXRegs_59_REG_2) : $signed(_GEN_1586); // @[\\src\\main\\scala\\GameLogic.scala 660:37 663:25]
  wire [9:0] _GEN_1595 = starCnt == 10'hf0 ? $signed(spriteYRegs_59_REG_2) : $signed(_GEN_1589); // @[\\src\\main\\scala\\GameLogic.scala 660:37 664:25]
  wire [10:0] _GEN_1596 = starCnt == 10'hf0 ? $signed(spriteXRegs_60_REG_2) : $signed(_GEN_1587); // @[\\src\\main\\scala\\GameLogic.scala 660:37 665:25]
  wire [9:0] _GEN_1597 = starCnt == 10'hf0 ? $signed(spriteYRegs_60_REG_2) : $signed(_GEN_1590); // @[\\src\\main\\scala\\GameLogic.scala 660:37 666:25]
  wire  _GEN_1598 = starCnt == 10'hf0 | _GEN_1579; // @[\\src\\main\\scala\\GameLogic.scala 660:37 667:35]
  wire  _GEN_1599 = starCnt == 10'hf0 | _GEN_1580; // @[\\src\\main\\scala\\GameLogic.scala 660:37 668:35]
  wire  _GEN_1600 = starCnt == 10'hf0 | _GEN_1581; // @[\\src\\main\\scala\\GameLogic.scala 660:37 669:35]
  wire  _GEN_1601 = starCnt == 10'hf0 | _GEN_1582; // @[\\src\\main\\scala\\GameLogic.scala 660:37 670:33]
  wire  _GEN_1602 = starCnt == 10'hf0 | _GEN_1583; // @[\\src\\main\\scala\\GameLogic.scala 660:37 671:33]
  wire  _GEN_1603 = starCnt == 10'hf0 | _GEN_1584; // @[\\src\\main\\scala\\GameLogic.scala 660:37 672:33]
  wire [9:0] _GEN_1604 = starCnt == 10'hf0 ? _starCnt_T_1 : _GEN_1591; // @[\\src\\main\\scala\\GameLogic.scala 660:37 673:17]
  wire  _GEN_1605 = starCnt == 10'hb4 ? 1'h0 : _GEN_1598; // @[\\src\\main\\scala\\GameLogic.scala 646:37 647:35]
  wire  _GEN_1606 = starCnt == 10'hb4 ? 1'h0 : _GEN_1599; // @[\\src\\main\\scala\\GameLogic.scala 646:37 648:35]
  wire  _GEN_1607 = starCnt == 10'hb4 ? 1'h0 : _GEN_1600; // @[\\src\\main\\scala\\GameLogic.scala 646:37 649:35]
  wire  _GEN_1608 = starCnt == 10'hb4 ? 1'h0 : _GEN_1601; // @[\\src\\main\\scala\\GameLogic.scala 646:37 650:33]
  wire  _GEN_1609 = starCnt == 10'hb4 ? 1'h0 : _GEN_1602; // @[\\src\\main\\scala\\GameLogic.scala 646:37 651:33]
  wire  _GEN_1610 = starCnt == 10'hb4 ? 1'h0 : _GEN_1603; // @[\\src\\main\\scala\\GameLogic.scala 646:37 652:33]
  wire [10:0] _GEN_1611 = starCnt == 10'hb4 ? $signed(_spriteXRegs_58_T_5) : $signed(_GEN_1592); // @[\\src\\main\\scala\\GameLogic.scala 646:37 653:25]
  wire [10:0] _GEN_1612 = starCnt == 10'hb4 ? $signed(_spriteXRegs_59_T_5) : $signed(_GEN_1594); // @[\\src\\main\\scala\\GameLogic.scala 646:37 654:25]
  wire [10:0] _GEN_1613 = starCnt == 10'hb4 ? $signed(_spriteXRegs_60_T_5) : $signed(_GEN_1596); // @[\\src\\main\\scala\\GameLogic.scala 646:37 655:25]
  wire [9:0] _GEN_1614 = starCnt == 10'hb4 ? $signed(_spriteYRegs_58_T_5) : $signed(_GEN_1593); // @[\\src\\main\\scala\\GameLogic.scala 646:37 656:25]
  wire [9:0] _GEN_1615 = starCnt == 10'hb4 ? $signed(_spriteYRegs_59_T_5) : $signed(_GEN_1595); // @[\\src\\main\\scala\\GameLogic.scala 646:37 657:25]
  wire [9:0] _GEN_1616 = starCnt == 10'hb4 ? $signed(_spriteYRegs_60_T_5) : $signed(_GEN_1597); // @[\\src\\main\\scala\\GameLogic.scala 646:37 658:25]
  wire [9:0] _GEN_1617 = starCnt == 10'hb4 ? _starCnt_T_1 : _GEN_1604; // @[\\src\\main\\scala\\GameLogic.scala 646:37 659:17]
  wire [10:0] _GEN_1618 = starCnt == 10'h78 ? $signed(spriteXRegs_58_REG_1) : $signed(_GEN_1611); // @[\\src\\main\\scala\\GameLogic.scala 632:37 633:25]
  wire [9:0] _GEN_1619 = starCnt == 10'h78 ? $signed(spriteYRegs_58_REG_1) : $signed(_GEN_1614); // @[\\src\\main\\scala\\GameLogic.scala 632:37 634:25]
  wire [10:0] _GEN_1620 = starCnt == 10'h78 ? $signed(spriteXRegs_59_REG_1) : $signed(_GEN_1612); // @[\\src\\main\\scala\\GameLogic.scala 632:37 635:25]
  wire [9:0] _GEN_1621 = starCnt == 10'h78 ? $signed(spriteYRegs_59_REG_1) : $signed(_GEN_1615); // @[\\src\\main\\scala\\GameLogic.scala 632:37 636:25]
  wire [10:0] _GEN_1622 = starCnt == 10'h78 ? $signed(spriteXRegs_60_REG_1) : $signed(_GEN_1613); // @[\\src\\main\\scala\\GameLogic.scala 632:37 637:25]
  wire [9:0] _GEN_1623 = starCnt == 10'h78 ? $signed(spriteYRegs_60_REG_1) : $signed(_GEN_1616); // @[\\src\\main\\scala\\GameLogic.scala 632:37 638:25]
  wire  _GEN_1624 = starCnt == 10'h78 | _GEN_1605; // @[\\src\\main\\scala\\GameLogic.scala 632:37 639:35]
  wire  _GEN_1625 = starCnt == 10'h78 | _GEN_1606; // @[\\src\\main\\scala\\GameLogic.scala 632:37 640:35]
  wire  _GEN_1626 = starCnt == 10'h78 | _GEN_1607; // @[\\src\\main\\scala\\GameLogic.scala 632:37 641:35]
  wire  _GEN_1627 = starCnt == 10'h78 | _GEN_1608; // @[\\src\\main\\scala\\GameLogic.scala 632:37 642:33]
  wire  _GEN_1628 = starCnt == 10'h78 | _GEN_1609; // @[\\src\\main\\scala\\GameLogic.scala 632:37 643:33]
  wire  _GEN_1629 = starCnt == 10'h78 | _GEN_1610; // @[\\src\\main\\scala\\GameLogic.scala 632:37 644:33]
  wire [9:0] _GEN_1630 = starCnt == 10'h78 ? _starCnt_T_1 : _GEN_1617; // @[\\src\\main\\scala\\GameLogic.scala 632:37 645:17]
  wire  _GEN_1631 = starCnt == 10'h3c ? 1'h0 : _GEN_1624; // @[\\src\\main\\scala\\GameLogic.scala 618:36 619:35]
  wire  _GEN_1632 = starCnt == 10'h3c ? 1'h0 : _GEN_1625; // @[\\src\\main\\scala\\GameLogic.scala 618:36 620:35]
  wire  _GEN_1633 = starCnt == 10'h3c ? 1'h0 : _GEN_1626; // @[\\src\\main\\scala\\GameLogic.scala 618:36 621:35]
  wire  _GEN_1634 = starCnt == 10'h3c ? 1'h0 : _GEN_1627; // @[\\src\\main\\scala\\GameLogic.scala 618:36 622:33]
  wire  _GEN_1635 = starCnt == 10'h3c ? 1'h0 : _GEN_1628; // @[\\src\\main\\scala\\GameLogic.scala 618:36 623:33]
  wire  _GEN_1636 = starCnt == 10'h3c ? 1'h0 : _GEN_1629; // @[\\src\\main\\scala\\GameLogic.scala 618:36 624:33]
  wire [10:0] _GEN_1637 = starCnt == 10'h3c ? $signed(_spriteXRegs_58_T_5) : $signed(_GEN_1618); // @[\\src\\main\\scala\\GameLogic.scala 618:36 625:25]
  wire [10:0] _GEN_1638 = starCnt == 10'h3c ? $signed(_spriteXRegs_59_T_5) : $signed(_GEN_1620); // @[\\src\\main\\scala\\GameLogic.scala 618:36 626:25]
  wire [10:0] _GEN_1639 = starCnt == 10'h3c ? $signed(_spriteXRegs_60_T_5) : $signed(_GEN_1622); // @[\\src\\main\\scala\\GameLogic.scala 618:36 627:25]
  wire [9:0] _GEN_1640 = starCnt == 10'h3c ? $signed(_spriteYRegs_58_T_5) : $signed(_GEN_1619); // @[\\src\\main\\scala\\GameLogic.scala 618:36 628:25]
  wire [9:0] _GEN_1641 = starCnt == 10'h3c ? $signed(_spriteYRegs_59_T_5) : $signed(_GEN_1621); // @[\\src\\main\\scala\\GameLogic.scala 618:36 629:25]
  wire [9:0] _GEN_1642 = starCnt == 10'h3c ? $signed(_spriteYRegs_60_T_5) : $signed(_GEN_1623); // @[\\src\\main\\scala\\GameLogic.scala 618:36 630:25]
  wire [9:0] _GEN_1643 = starCnt == 10'h3c ? _starCnt_T_1 : _GEN_1630; // @[\\src\\main\\scala\\GameLogic.scala 618:36 631:17]
  wire  _GEN_1650 = starCnt == 10'h0 | _GEN_1631; // @[\\src\\main\\scala\\GameLogic.scala 604:29 611:35]
  wire  _GEN_1651 = starCnt == 10'h0 | _GEN_1632; // @[\\src\\main\\scala\\GameLogic.scala 604:29 612:35]
  wire  _GEN_1652 = starCnt == 10'h0 | _GEN_1633; // @[\\src\\main\\scala\\GameLogic.scala 604:29 613:35]
  wire  _GEN_1653 = starCnt == 10'h0 | _GEN_1634; // @[\\src\\main\\scala\\GameLogic.scala 604:29 614:33]
  wire  _GEN_1654 = starCnt == 10'h0 | _GEN_1635; // @[\\src\\main\\scala\\GameLogic.scala 604:29 615:33]
  wire  _GEN_1655 = starCnt == 10'h0 | _GEN_1636; // @[\\src\\main\\scala\\GameLogic.scala 604:29 616:33]
  wire  _T_815 = $signed(spriteYRegs_3) > 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 712:81]
  wire  _T_817 = $signed(spriteYRegs_3) < 10'sh14c; // @[\\src\\main\\scala\\GameLogic.scala 712:107]
  wire  _T_818 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c; // @[\\src\\main\\scala\\GameLogic.scala 712:89]
  wire [1:0] _GEN_1658 = io_btnC ? 2'h1 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 715:25 716:20 219:23]
  wire [2:0] _GEN_1659 = io_btnC ? 3'h3 : 3'h4; // @[\\src\\main\\scala\\GameLogic.scala 715:25 717:22 719:22]
  wire  _T_825 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817; // @[\\src\\main\\scala\\GameLogic.scala 721:95]
  wire [1:0] _GEN_1660 = io_btnC ? 2'h2 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 724:25 725:20 219:23]
  wire  _T_832 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_815 & _T_817; // @[\\src\\main\\scala\\GameLogic.scala 730:95]
  wire [1:0] _GEN_1661 = io_btnC ? 2'h3 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 733:25 734:20 219:23]
  wire  _GEN_1662 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_815 & _T_817 ? 1'h0 : 1'h1
    ; // @[\\src\\main\\scala\\GameLogic.scala 730:122 709:31 731:33]
  wire [1:0] _GEN_1664 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_815 & _T_817 ?
    _GEN_1661 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 730:122 219:23]
  wire [2:0] _GEN_1665 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_815 & _T_817 ?
    _GEN_1659 : 3'h4; // @[\\src\\main\\scala\\GameLogic.scala 730:122 740:20]
  wire  _GEN_1666 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 ? 1'h0 : 1'h1
    ; // @[\\src\\main\\scala\\GameLogic.scala 721:122 707:30 722:32]
  wire [1:0] _GEN_1668 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 ?
    _GEN_1660 : _GEN_1664; // @[\\src\\main\\scala\\GameLogic.scala 721:122]
  wire [2:0] _GEN_1669 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 ?
    _GEN_1659 : _GEN_1665; // @[\\src\\main\\scala\\GameLogic.scala 721:122]
  wire  _GEN_1670 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 | _GEN_1662; // @[\\src\\main\\scala\\GameLogic.scala 721:122 709:31]
  wire  _GEN_1671 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 ? 1'h0 :
    _T_832; // @[\\src\\main\\scala\\GameLogic.scala 721:122 710:31]
  wire  _GEN_1672 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 712:116 705:30 713:32]
  wire [1:0] _GEN_1674 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3)
     > 10'sh12c & $signed(spriteYRegs_3) < 10'sh14c ? _GEN_1658 : _GEN_1668; // @[\\src\\main\\scala\\GameLogic.scala 712:116]
  wire [2:0] _GEN_1675 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3)
     > 10'sh12c & $signed(spriteYRegs_3) < 10'sh14c ? _GEN_1659 : _GEN_1669; // @[\\src\\main\\scala\\GameLogic.scala 712:116]
  wire  _GEN_1676 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c | _GEN_1666; // @[\\src\\main\\scala\\GameLogic.scala 712:116 707:30]
  wire  _GEN_1677 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c ? 1'h0 : _T_825; // @[\\src\\main\\scala\\GameLogic.scala 712:116 708:31]
  wire  _GEN_1678 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c | _GEN_1670; // @[\\src\\main\\scala\\GameLogic.scala 712:116 709:31]
  wire  _GEN_1679 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c ? 1'h0 : _GEN_1671; // @[\\src\\main\\scala\\GameLogic.scala 712:116 710:31]
  wire [2:0] _GEN_1680 = _T ? 3'h4 : _GEN_1675; // @[\\src\\main\\scala\\GameLogic.scala 700:28 701:18]
  wire  _GEN_1681 = _T ? spriteVisibleRegs_3 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 700:28 125:34 704:30]
  wire  _GEN_1682 = _T ? spriteVisibleRegs_7 : _GEN_1672; // @[\\src\\main\\scala\\GameLogic.scala 700:28 125:34]
  wire  _GEN_1683 = _T ? spriteVisibleRegs_8 : _T_818; // @[\\src\\main\\scala\\GameLogic.scala 700:28 125:34]
  wire  _GEN_1684 = _T ? spriteVisibleRegs_9 : _GEN_1676; // @[\\src\\main\\scala\\GameLogic.scala 700:28 125:34]
  wire  _GEN_1685 = _T ? spriteVisibleRegs_10 : _GEN_1677; // @[\\src\\main\\scala\\GameLogic.scala 700:28 125:34]
  wire  _GEN_1686 = _T ? spriteVisibleRegs_11 : _GEN_1678; // @[\\src\\main\\scala\\GameLogic.scala 700:28 125:34]
  wire  _GEN_1687 = _T ? spriteVisibleRegs_12 : _GEN_1679; // @[\\src\\main\\scala\\GameLogic.scala 700:28 125:34]
  wire [1:0] _GEN_1688 = _T ? lvlReg : _GEN_1674; // @[\\src\\main\\scala\\GameLogic.scala 219:23 700:28]
  wire [9:0] _GEN_1689 = _T_83 ? 10'h280 : viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 768:34 769:21 209:28]
  wire [8:0] _GEN_1690 = _T_83 ? 9'h1e0 : viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 768:34 770:21 210:28]
  wire [9:0] _GEN_1691 = _T_76 ? 10'h0 : _GEN_1689; // @[\\src\\main\\scala\\GameLogic.scala 765:34 766:21]
  wire [8:0] _GEN_1692 = _T_76 ? 9'h1e0 : _GEN_1690; // @[\\src\\main\\scala\\GameLogic.scala 765:34 767:21]
  wire [9:0] _GEN_1693 = _T_69 ? 10'h280 : _GEN_1691; // @[\\src\\main\\scala\\GameLogic.scala 762:28 763:21]
  wire [8:0] _GEN_1694 = _T_69 ? 9'h0 : _GEN_1692; // @[\\src\\main\\scala\\GameLogic.scala 762:28 764:21]
  wire [9:0] _spriteYRegs_14_T_2 = $signed(spriteYRegs_14) + 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 780:48]
  wire [9:0] _GEN_1695 = $signed(spriteYRegs_14) < 10'sh1c0 ? $signed(_spriteYRegs_14_T_2) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 779:48 780:29]
  wire [9:0] _spriteYRegs_14_T_5 = $signed(spriteYRegs_14) - 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 784:48]
  wire [9:0] _GEN_1696 = $signed(spriteYRegs_14) > 10'sh20 ? $signed(_spriteYRegs_14_T_5) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 783:40 784:29]
  wire [9:0] _GEN_1697 = io_btnU ? $signed(_GEN_1696) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 782:29]
  wire [9:0] _GEN_1698 = io_btnD ? $signed(_GEN_1695) : $signed(_GEN_1697); // @[\\src\\main\\scala\\GameLogic.scala 778:23]
  wire [9:0] _spriteYRegs_3_T_2 = $signed(spriteYRegs_3) + 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 323:58]
  wire [9:0] _GEN_1699 = $signed(spriteYRegs_3) < 10'sh1c0 ? $signed(_spriteYRegs_3_T_2) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 322:51 323:32]
  wire [9:0] _spriteYRegs_3_T_5 = $signed(spriteYRegs_3) - 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 327:58]
  wire [9:0] _GEN_1700 = $signed(spriteYRegs_3) > 10'sh20 ? $signed(_spriteYRegs_3_T_5) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 326:43 327:32]
  wire [9:0] _GEN_1701 = io_btnU ? $signed(_GEN_1700) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 325:25]
  wire [9:0] _GEN_1702 = io_btnD ? $signed(_GEN_1699) : $signed(_GEN_1701); // @[\\src\\main\\scala\\GameLogic.scala 321:19]
  wire [10:0] _spriteXRegs_3_T_2 = $signed(spriteXRegs_3) + 11'sh2; // @[\\src\\main\\scala\\GameLogic.scala 332:58]
  wire [10:0] _GEN_1703 = $signed(spriteXRegs_3) < 11'sh260 ? $signed(_spriteXRegs_3_T_2) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 331:51 332:32]
  wire [10:0] _spriteXRegs_3_T_5 = $signed(spriteXRegs_3) - 11'sh2; // @[\\src\\main\\scala\\GameLogic.scala 336:58]
  wire [10:0] _GEN_1704 = $signed(spriteXRegs_3) > 11'sh20 ? $signed(_spriteXRegs_3_T_5) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 335:43 336:32]
  wire [10:0] _GEN_1705 = io_btnL ? $signed(_GEN_1704) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 334:25]
  wire [10:0] _GEN_1706 = io_btnR ? $signed(_GEN_1703) : $signed(_GEN_1705); // @[\\src\\main\\scala\\GameLogic.scala 330:19]
  wire [9:0] _GEN_1707 = _T ? $signed(_GEN_1698) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 777:28]
  wire [9:0] _GEN_1708 = _T ? $signed(_GEN_1) : $signed(_GEN_1702); // @[\\src\\main\\scala\\GameLogic.scala 777:28]
  wire [10:0] _GEN_1709 = _T ? $signed(_GEN_0) : $signed(_GEN_1706); // @[\\src\\main\\scala\\GameLogic.scala 777:28]
  wire [2:0] _GEN_1710 = _T_5 ? 3'h6 : 3'h5; // @[\\src\\main\\scala\\GameLogic.scala 792:30 793:18 795:18]
  wire [10:0] _cursorOnReturn_T_2 = $signed(spriteXRegs_3) + 11'sh1c; // @[\\src\\main\\scala\\GameLogic.scala 810:44]
  wire [9:0] _cursorOnReturn_T_11 = $signed(spriteYRegs_3) + 10'sh7; // @[\\src\\main\\scala\\GameLogic.scala 811:25]
  wire  _cursorOnReturn_T_12 = $signed(_cursorOnReturn_T_11) >= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 811:32]
  wire  _cursorOnReturn_T_13 = $signed(_cursorOnReturn_T_2) >= 11'sh110 & $signed(_cursorOnReturn_T_2) <= 11'sh170 &
    _cursorOnReturn_T_12; // @[\\src\\main\\scala\\GameLogic.scala 810:97]
  wire  cursorOnReturn = _cursorOnReturn_T_13 & $signed(_cursorOnReturn_T_11) <= 10'sh124; // @[\\src\\main\\scala\\GameLogic.scala 811:41]
  wire  _spriteVisibleRegs_52_T = ~cursorOnReturn; // @[\\src\\main\\scala\\GameLogic.scala 813:32]
  wire  _GEN_1719 = cursorOnReturn & io_btnC | gameOverReturnPressed; // @[\\src\\main\\scala\\GameLogic.scala 825:39 826:31 237:38]
  wire [2:0] _GEN_1722 = 3'h5 == stateReg ? 3'h0 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 346:20 835:16 113:25]
  wire  _GEN_1723 = 3'h6 == stateReg ? 1'h0 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 346:20 800:29 125:34]
  wire  _GEN_1724 = 3'h6 == stateReg | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 346:20 803:29 125:34]
  wire  _GEN_1725 = 3'h6 == stateReg | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 346:20 804:29 125:34]
  wire  _GEN_1726 = 3'h6 == stateReg | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 346:20 805:29 125:34]
  wire  _GEN_1727 = 3'h6 == stateReg | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 346:20 806:29 125:34]
  wire  _GEN_1728 = 3'h6 == stateReg | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 346:20 807:29 125:34]
  wire  _GEN_1729 = 3'h6 == stateReg | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 346:20 808:29 125:34]
  wire  _GEN_1730 = 3'h6 == stateReg ? ~cursorOnReturn : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 346:20 813:29 125:34]
  wire  _GEN_1731 = 3'h6 == stateReg ? _spriteVisibleRegs_52_T : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 346:20 814:29 125:34]
  wire  _GEN_1732 = 3'h6 == stateReg ? _spriteVisibleRegs_52_T : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 346:20 815:29 125:34]
  wire  _GEN_1733 = 3'h6 == stateReg ? cursorOnReturn : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 346:20 816:29 125:34]
  wire  _GEN_1734 = 3'h6 == stateReg ? cursorOnReturn : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 346:20 817:29 125:34]
  wire  _GEN_1735 = 3'h6 == stateReg ? cursorOnReturn : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 346:20 818:29 125:34]
  wire  _GEN_1736 = 3'h6 == stateReg | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 346:20 821:28 125:34]
  wire [9:0] _GEN_1737 = 3'h6 == stateReg ? $signed(_GEN_1702) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [10:0] _GEN_1738 = 3'h6 == stateReg ? $signed(_GEN_1706) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1739 = 3'h6 == stateReg ? _GEN_1719 : gameOverReturnPressed; // @[\\src\\main\\scala\\GameLogic.scala 346:20 237:38]
  wire [2:0] _GEN_1741 = 3'h6 == stateReg ? 3'h5 : _GEN_1722; // @[\\src\\main\\scala\\GameLogic.scala 346:20 831:16]
  wire  _GEN_1742 = 3'h6 == stateReg ? 1'h0 : 3'h5 == stateReg; // @[\\src\\main\\scala\\GameLogic.scala 346:20 100:22]
  wire [9:0] _GEN_1743 = 3'h4 == stateReg ? $signed(_GEN_1707) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [9:0] _GEN_1744 = 3'h4 == stateReg ? $signed(_GEN_1708) : $signed(_GEN_1737); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [10:0] _GEN_1745 = 3'h4 == stateReg ? $signed(_GEN_1709) : $signed(_GEN_1738); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [2:0] _GEN_1746 = 3'h4 == stateReg ? _GEN_1710 : _GEN_1741; // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1747 = 3'h4 == stateReg ? spriteVisibleRegs_14 : _GEN_1723; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1748 = 3'h4 == stateReg ? spriteVisibleRegs_46 : _GEN_1724; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1749 = 3'h4 == stateReg ? spriteVisibleRegs_47 : _GEN_1725; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1750 = 3'h4 == stateReg ? spriteVisibleRegs_48 : _GEN_1726; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1751 = 3'h4 == stateReg ? spriteVisibleRegs_49 : _GEN_1727; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1752 = 3'h4 == stateReg ? spriteVisibleRegs_50 : _GEN_1728; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1753 = 3'h4 == stateReg ? spriteVisibleRegs_51 : _GEN_1729; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1754 = 3'h4 == stateReg ? spriteVisibleRegs_52 : _GEN_1730; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1755 = 3'h4 == stateReg ? spriteVisibleRegs_53 : _GEN_1731; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1756 = 3'h4 == stateReg ? spriteVisibleRegs_54 : _GEN_1732; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1757 = 3'h4 == stateReg ? spriteVisibleRegs_55 : _GEN_1733; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1758 = 3'h4 == stateReg ? spriteVisibleRegs_56 : _GEN_1734; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1759 = 3'h4 == stateReg ? spriteVisibleRegs_57 : _GEN_1735; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1760 = 3'h4 == stateReg ? spriteVisibleRegs_3 : _GEN_1736; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1761 = 3'h4 == stateReg ? gameOverReturnPressed : _GEN_1739; // @[\\src\\main\\scala\\GameLogic.scala 346:20 237:38]
  wire  _GEN_1763 = 3'h4 == stateReg ? 1'h0 : _GEN_1742; // @[\\src\\main\\scala\\GameLogic.scala 346:20 100:22]
  wire [5:0] _GEN_1764 = 3'h3 == stateReg ? 6'h0 : nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 346:20 746:25 244:34]
  wire [7:0] _GEN_1765 = 3'h3 == stateReg ? 8'h0 : spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 346:20 747:25 243:34]
  wire [10:0] _GEN_1766 = 3'h3 == stateReg ? $signed(11'sh260) : $signed(_GEN_16); // @[\\src\\main\\scala\\GameLogic.scala 346:20 749:23]
  wire [9:0] _GEN_1767 = 3'h3 == stateReg ? $signed(10'sh140) : $signed(_GEN_1743); // @[\\src\\main\\scala\\GameLogic.scala 346:20 750:23]
  wire  _GEN_1768 = 3'h3 == stateReg ? 1'h0 : _GEN_1760; // @[\\src\\main\\scala\\GameLogic.scala 346:20 751:28]
  wire  _GEN_1769 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 346:20 752:28 125:34]
  wire  _GEN_1770 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 346:20 753:28 125:34]
  wire  _GEN_1771 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 346:20 754:28 125:34]
  wire  _GEN_1772 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 346:20 755:29 125:34]
  wire  _GEN_1773 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 346:20 756:29 125:34]
  wire  _GEN_1774 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 346:20 757:29 125:34]
  wire  _GEN_1775 = 3'h3 == stateReg | _GEN_1747; // @[\\src\\main\\scala\\GameLogic.scala 346:20 758:29]
  wire  _GEN_1776 = 3'h3 == stateReg | _GEN_195; // @[\\src\\main\\scala\\GameLogic.scala 346:20 759:29]
  wire  _GEN_1777 = 3'h3 == stateReg | _GEN_196; // @[\\src\\main\\scala\\GameLogic.scala 346:20 760:29]
  wire  _GEN_1778 = 3'h3 == stateReg | _GEN_197; // @[\\src\\main\\scala\\GameLogic.scala 346:20 761:29]
  wire [9:0] _GEN_1779 = 3'h3 == stateReg ? _GEN_1693 : viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 346:20 209:28]
  wire [8:0] _GEN_1780 = 3'h3 == stateReg ? _GEN_1694 : viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 346:20 210:28]
  wire [2:0] _GEN_1781 = 3'h3 == stateReg ? 3'h4 : _GEN_1746; // @[\\src\\main\\scala\\GameLogic.scala 346:20 772:16]
  wire [9:0] _GEN_1782 = 3'h3 == stateReg ? $signed(_GEN_1) : $signed(_GEN_1744); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [10:0] _GEN_1783 = 3'h3 == stateReg ? $signed(_GEN_0) : $signed(_GEN_1745); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1784 = 3'h3 == stateReg ? spriteVisibleRegs_46 : _GEN_1748; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1785 = 3'h3 == stateReg ? spriteVisibleRegs_47 : _GEN_1749; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1786 = 3'h3 == stateReg ? spriteVisibleRegs_48 : _GEN_1750; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1787 = 3'h3 == stateReg ? spriteVisibleRegs_49 : _GEN_1751; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1788 = 3'h3 == stateReg ? spriteVisibleRegs_50 : _GEN_1752; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1789 = 3'h3 == stateReg ? spriteVisibleRegs_51 : _GEN_1753; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1790 = 3'h3 == stateReg ? spriteVisibleRegs_52 : _GEN_1754; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1791 = 3'h3 == stateReg ? spriteVisibleRegs_53 : _GEN_1755; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1792 = 3'h3 == stateReg ? spriteVisibleRegs_54 : _GEN_1756; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1793 = 3'h3 == stateReg ? spriteVisibleRegs_55 : _GEN_1757; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1794 = 3'h3 == stateReg ? spriteVisibleRegs_56 : _GEN_1758; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1795 = 3'h3 == stateReg ? spriteVisibleRegs_57 : _GEN_1759; // @[\\src\\main\\scala\\GameLogic.scala 346:20 125:34]
  wire  _GEN_1796 = 3'h3 == stateReg ? gameOverReturnPressed : _GEN_1761; // @[\\src\\main\\scala\\GameLogic.scala 346:20 237:38]
  wire  _GEN_1798 = 3'h3 == stateReg ? 1'h0 : _GEN_1763; // @[\\src\\main\\scala\\GameLogic.scala 346:20 100:22]
  wire  _GEN_1834 = 3'h2 == stateReg ? 1'h0 : _GEN_1798; // @[\\src\\main\\scala\\GameLogic.scala 346:20 100:22]
  wire [26:0] _GEN_1837 = 3'h1 == stateReg ? $signed(_GEN_471) : $signed({{16{_GEN_18[10]}},_GEN_18}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1840 = 3'h1 == stateReg ? _GEN_474 : spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1842 = 3'h1 == stateReg ? $signed(_GEN_476) : $signed({{16{_GEN_20[10]}},_GEN_20}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1845 = 3'h1 == stateReg ? _GEN_479 : spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1847 = 3'h1 == stateReg ? $signed(_GEN_481) : $signed({{16{_GEN_22[10]}},_GEN_22}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1850 = 3'h1 == stateReg ? _GEN_484 : spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1852 = 3'h1 == stateReg ? $signed(_GEN_486) : $signed({{16{_GEN_24[10]}},_GEN_24}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1855 = 3'h1 == stateReg ? _GEN_489 : spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1857 = 3'h1 == stateReg ? $signed(_GEN_491) : $signed({{16{_GEN_26[10]}},_GEN_26}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1860 = 3'h1 == stateReg ? _GEN_494 : spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1862 = 3'h1 == stateReg ? $signed(_GEN_496) : $signed({{16{_GEN_28[10]}},_GEN_28}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1865 = 3'h1 == stateReg ? _GEN_499 : spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1867 = 3'h1 == stateReg ? $signed(_GEN_501) : $signed({{16{_GEN_30[10]}},_GEN_30}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1870 = 3'h1 == stateReg ? _GEN_504 : spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1872 = 3'h1 == stateReg ? $signed(_GEN_506) : $signed({{16{_GEN_32[10]}},_GEN_32}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1875 = 3'h1 == stateReg ? _GEN_509 : spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1877 = 3'h1 == stateReg ? $signed(_GEN_511) : $signed({{16{_GEN_34[10]}},_GEN_34}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1880 = 3'h1 == stateReg ? _GEN_514 : spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1882 = 3'h1 == stateReg ? $signed(_GEN_516) : $signed({{16{_GEN_36[10]}},_GEN_36}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_1885 = 3'h1 == stateReg ? _GEN_519 : spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  wire [26:0] _GEN_1887 = 3'h1 == stateReg ? $signed(_GEN_521) : $signed({{16{_GEN_38[10]}},_GEN_38}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1891 = 3'h1 == stateReg ? $signed(_GEN_525) : $signed({{16{_GEN_40[10]}},_GEN_40}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1895 = 3'h1 == stateReg ? $signed(_GEN_529) : $signed({{16{_GEN_42[10]}},_GEN_42}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1899 = 3'h1 == stateReg ? $signed(_GEN_533) : $signed({{16{_GEN_44[10]}},_GEN_44}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1903 = 3'h1 == stateReg ? $signed(_GEN_537) : $signed({{16{_GEN_46[10]}},_GEN_46}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1907 = 3'h1 == stateReg ? $signed(_GEN_541) : $signed({{16{_GEN_48[10]}},_GEN_48}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1911 = 3'h1 == stateReg ? $signed(_GEN_545) : $signed({{16{_GEN_50[10]}},_GEN_50}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1915 = 3'h1 == stateReg ? $signed(_GEN_549) : $signed({{16{_GEN_52[10]}},_GEN_52}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1919 = 3'h1 == stateReg ? $signed(_GEN_553) : $signed({{16{_GEN_54[10]}},_GEN_54}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1923 = 3'h1 == stateReg ? $signed(_GEN_557) : $signed({{16{_GEN_56[10]}},_GEN_56}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1927 = 3'h1 == stateReg ? $signed(_GEN_561) : $signed({{16{_GEN_58[10]}},_GEN_58}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1931 = 3'h1 == stateReg ? $signed(_GEN_565) : $signed({{16{_GEN_60[10]}},_GEN_60}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1935 = 3'h1 == stateReg ? $signed(_GEN_569) : $signed({{16{_GEN_62[10]}},_GEN_62}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1939 = 3'h1 == stateReg ? $signed(_GEN_573) : $signed({{16{_GEN_64[10]}},_GEN_64}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1943 = 3'h1 == stateReg ? $signed(_GEN_577) : $signed({{16{_GEN_66[10]}},_GEN_66}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1947 = 3'h1 == stateReg ? $signed(_GEN_581) : $signed({{16{_GEN_68[10]}},_GEN_68}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1951 = 3'h1 == stateReg ? $signed(_GEN_585) : $signed({{16{_GEN_70[10]}},_GEN_70}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1955 = 3'h1 == stateReg ? $signed(_GEN_589) : $signed({{16{_GEN_72[10]}},_GEN_72}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1959 = 3'h1 == stateReg ? $signed(_GEN_593) : $signed({{16{_GEN_74[10]}},_GEN_74}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_1963 = 3'h1 == stateReg ? $signed(_GEN_597) : $signed({{16{_GEN_76[10]}},_GEN_76}); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire  _GEN_2100 = 3'h1 == stateReg ? 1'h0 : _GEN_1834; // @[\\src\\main\\scala\\GameLogic.scala 346:20 100:22]
  wire  _GEN_2112 = 3'h0 == stateReg ? _GEN_268 : _GEN_186; // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2160 = 3'h0 == stateReg ? $signed({{16{_GEN_18[10]}},_GEN_18}) : $signed(_GEN_1837); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2165 = 3'h0 == stateReg ? $signed({{16{_GEN_20[10]}},_GEN_20}) : $signed(_GEN_1842); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2170 = 3'h0 == stateReg ? $signed({{16{_GEN_22[10]}},_GEN_22}) : $signed(_GEN_1847); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2175 = 3'h0 == stateReg ? $signed({{16{_GEN_24[10]}},_GEN_24}) : $signed(_GEN_1852); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2180 = 3'h0 == stateReg ? $signed({{16{_GEN_26[10]}},_GEN_26}) : $signed(_GEN_1857); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2185 = 3'h0 == stateReg ? $signed({{16{_GEN_28[10]}},_GEN_28}) : $signed(_GEN_1862); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2190 = 3'h0 == stateReg ? $signed({{16{_GEN_30[10]}},_GEN_30}) : $signed(_GEN_1867); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2195 = 3'h0 == stateReg ? $signed({{16{_GEN_32[10]}},_GEN_32}) : $signed(_GEN_1872); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2200 = 3'h0 == stateReg ? $signed({{16{_GEN_34[10]}},_GEN_34}) : $signed(_GEN_1877); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2205 = 3'h0 == stateReg ? $signed({{16{_GEN_36[10]}},_GEN_36}) : $signed(_GEN_1882); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2210 = 3'h0 == stateReg ? $signed({{16{_GEN_38[10]}},_GEN_38}) : $signed(_GEN_1887); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2214 = 3'h0 == stateReg ? $signed({{16{_GEN_40[10]}},_GEN_40}) : $signed(_GEN_1891); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2218 = 3'h0 == stateReg ? $signed({{16{_GEN_42[10]}},_GEN_42}) : $signed(_GEN_1895); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2222 = 3'h0 == stateReg ? $signed({{16{_GEN_44[10]}},_GEN_44}) : $signed(_GEN_1899); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2226 = 3'h0 == stateReg ? $signed({{16{_GEN_46[10]}},_GEN_46}) : $signed(_GEN_1903); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2230 = 3'h0 == stateReg ? $signed({{16{_GEN_48[10]}},_GEN_48}) : $signed(_GEN_1907); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2234 = 3'h0 == stateReg ? $signed({{16{_GEN_50[10]}},_GEN_50}) : $signed(_GEN_1911); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2238 = 3'h0 == stateReg ? $signed({{16{_GEN_52[10]}},_GEN_52}) : $signed(_GEN_1915); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2242 = 3'h0 == stateReg ? $signed({{16{_GEN_54[10]}},_GEN_54}) : $signed(_GEN_1919); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2246 = 3'h0 == stateReg ? $signed({{16{_GEN_56[10]}},_GEN_56}) : $signed(_GEN_1923); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2250 = 3'h0 == stateReg ? $signed({{16{_GEN_58[10]}},_GEN_58}) : $signed(_GEN_1927); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2254 = 3'h0 == stateReg ? $signed({{16{_GEN_60[10]}},_GEN_60}) : $signed(_GEN_1931); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2258 = 3'h0 == stateReg ? $signed({{16{_GEN_62[10]}},_GEN_62}) : $signed(_GEN_1935); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2262 = 3'h0 == stateReg ? $signed({{16{_GEN_64[10]}},_GEN_64}) : $signed(_GEN_1939); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2266 = 3'h0 == stateReg ? $signed({{16{_GEN_66[10]}},_GEN_66}) : $signed(_GEN_1943); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2270 = 3'h0 == stateReg ? $signed({{16{_GEN_68[10]}},_GEN_68}) : $signed(_GEN_1947); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2274 = 3'h0 == stateReg ? $signed({{16{_GEN_70[10]}},_GEN_70}) : $signed(_GEN_1951); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2278 = 3'h0 == stateReg ? $signed({{16{_GEN_72[10]}},_GEN_72}) : $signed(_GEN_1955); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2282 = 3'h0 == stateReg ? $signed({{16{_GEN_74[10]}},_GEN_74}) : $signed(_GEN_1959); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2286 = 3'h0 == stateReg ? $signed({{16{_GEN_76[10]}},_GEN_76}) : $signed(_GEN_1963); // @[\\src\\main\\scala\\GameLogic.scala 346:20]
  wire [26:0] _GEN_2775 = reset ? $signed(27'sh0) : $signed(_GEN_2160); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2777 = reset ? $signed(27'sh0) : $signed(_GEN_2165); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2779 = reset ? $signed(27'sh0) : $signed(_GEN_2170); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2781 = reset ? $signed(27'sh0) : $signed(_GEN_2175); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2783 = reset ? $signed(27'sh0) : $signed(_GEN_2180); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2785 = reset ? $signed(27'sh0) : $signed(_GEN_2185); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2787 = reset ? $signed(27'sh0) : $signed(_GEN_2190); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2789 = reset ? $signed(27'sh0) : $signed(_GEN_2195); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2791 = reset ? $signed(27'sh0) : $signed(_GEN_2200); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2793 = reset ? $signed(27'sh0) : $signed(_GEN_2205); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2795 = reset ? $signed(27'sh0) : $signed(_GEN_2210); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2797 = reset ? $signed(27'sh0) : $signed(_GEN_2214); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2799 = reset ? $signed(27'sh0) : $signed(_GEN_2218); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2801 = reset ? $signed(27'sh0) : $signed(_GEN_2222); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2803 = reset ? $signed(27'sh0) : $signed(_GEN_2226); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2805 = reset ? $signed(27'sh0) : $signed(_GEN_2230); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2807 = reset ? $signed(27'sh0) : $signed(_GEN_2234); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2809 = reset ? $signed(27'sh0) : $signed(_GEN_2238); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2811 = reset ? $signed(27'sh0) : $signed(_GEN_2242); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2813 = reset ? $signed(27'sh0) : $signed(_GEN_2246); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2815 = reset ? $signed(27'sh0) : $signed(_GEN_2250); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2817 = reset ? $signed(27'sh0) : $signed(_GEN_2254); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2819 = reset ? $signed(27'sh0) : $signed(_GEN_2258); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2821 = reset ? $signed(27'sh0) : $signed(_GEN_2262); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2823 = reset ? $signed(27'sh0) : $signed(_GEN_2266); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2825 = reset ? $signed(27'sh0) : $signed(_GEN_2270); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2827 = reset ? $signed(27'sh0) : $signed(_GEN_2274); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2829 = reset ? $signed(27'sh0) : $signed(_GEN_2278); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2831 = reset ? $signed(27'sh0) : $signed(_GEN_2282); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2833 = reset ? $signed(27'sh0) : $signed(_GEN_2286); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  Difficulty difficulty ( // @[\\src\\main\\scala\\GameLogic.scala 217:26]
    .clock(difficulty_clock),
    .reset(difficulty_reset),
    .io_level(difficulty_io_level),
    .io_speed(difficulty_io_speed),
    .io_resetSpeed(difficulty_io_resetSpeed)
  );
  LFSR lfsr ( // @[\\src\\main\\scala\\GameLogic.scala 259:20]
    .clock(lfsr_clock),
    .reset(lfsr_reset),
    .io_out_0(lfsr_io_out_0),
    .io_out_1(lfsr_io_out_1),
    .io_out_2(lfsr_io_out_2),
    .io_out_3(lfsr_io_out_3),
    .io_out_4(lfsr_io_out_4),
    .io_out_5(lfsr_io_out_5),
    .io_out_6(lfsr_io_out_6),
    .io_out_7(lfsr_io_out_7),
    .io_out_8(lfsr_io_out_8),
    .io_out_9(lfsr_io_out_9),
    .io_out_10(lfsr_io_out_10),
    .io_out_11(lfsr_io_out_11),
    .io_out_12(lfsr_io_out_12),
    .io_out_13(lfsr_io_out_13),
    .io_out_14(lfsr_io_out_14),
    .io_out_15(lfsr_io_out_15),
    .io_out_16(lfsr_io_out_16),
    .io_out_17(lfsr_io_out_17),
    .io_out_18(lfsr_io_out_18),
    .io_out_19(lfsr_io_out_19),
    .io_out_20(lfsr_io_out_20),
    .io_out_21(lfsr_io_out_21),
    .io_out_22(lfsr_io_out_22),
    .io_out_23(lfsr_io_out_23),
    .io_out_24(lfsr_io_out_24),
    .io_out_25(lfsr_io_out_25),
    .io_out_26(lfsr_io_out_26),
    .io_out_27(lfsr_io_out_27),
    .io_out_28(lfsr_io_out_28),
    .io_out_29(lfsr_io_out_29)
  );
  assign io_spriteXPosition_3 = spriteXRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_7 = spriteXRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_8 = spriteXRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_9 = spriteXRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_10 = spriteXRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_11 = spriteXRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_12 = spriteXRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_13 = spriteXRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_14 = spriteXRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_16 = spriteXRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_17 = spriteXRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_18 = spriteXRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_19 = spriteXRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_20 = spriteXRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_21 = spriteXRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_22 = spriteXRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_23 = spriteXRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_24 = spriteXRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_25 = spriteXRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_26 = spriteXRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_27 = spriteXRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_28 = spriteXRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_29 = spriteXRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_30 = spriteXRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_31 = spriteXRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_32 = spriteXRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_33 = spriteXRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_34 = spriteXRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_35 = spriteXRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_36 = spriteXRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_37 = spriteXRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_38 = spriteXRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_39 = spriteXRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_40 = spriteXRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_41 = spriteXRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_42 = spriteXRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_43 = spriteXRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_44 = spriteXRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_45 = spriteXRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_46 = spriteXRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_47 = spriteXRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_48 = spriteXRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_49 = spriteXRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_50 = spriteXRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_51 = spriteXRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_52 = spriteXRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_53 = spriteXRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_54 = spriteXRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_55 = spriteXRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_56 = spriteXRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_57 = spriteXRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_58 = spriteXRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_59 = spriteXRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_60 = spriteXRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_61 = spriteXRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_62 = spriteXRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteXPosition_63 = spriteXRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 188:27]
  assign io_spriteYPosition_3 = spriteYRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_7 = spriteYRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_8 = spriteYRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_9 = spriteYRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_10 = spriteYRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_11 = spriteYRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_12 = spriteYRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_13 = spriteYRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_14 = spriteYRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_16 = spriteYRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_17 = spriteYRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_18 = spriteYRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_19 = spriteYRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_20 = spriteYRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_21 = spriteYRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_22 = spriteYRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_23 = spriteYRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_24 = spriteYRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_25 = spriteYRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_26 = spriteYRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_27 = spriteYRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_28 = spriteYRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_29 = spriteYRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_30 = spriteYRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_31 = spriteYRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_32 = spriteYRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_33 = spriteYRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_34 = spriteYRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_35 = spriteYRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_36 = spriteYRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_37 = spriteYRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_38 = spriteYRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_39 = spriteYRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_40 = spriteYRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_41 = spriteYRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_42 = spriteYRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_43 = spriteYRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_44 = spriteYRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_45 = spriteYRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_46 = spriteYRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_47 = spriteYRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_48 = spriteYRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_49 = spriteYRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_50 = spriteYRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_51 = spriteYRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_52 = spriteYRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_53 = spriteYRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_54 = spriteYRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_55 = spriteYRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_56 = spriteYRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_57 = spriteYRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_58 = spriteYRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_59 = spriteYRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_60 = spriteYRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_61 = spriteYRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_62 = spriteYRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteYPosition_63 = spriteYRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 189:27]
  assign io_spriteVisible_3 = spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_4 = spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_5 = spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_6 = spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_7 = spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_8 = spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_9 = spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_10 = spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_11 = spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_12 = spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_13 = spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_14 = spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_15 = spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_16 = spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_17 = spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_18 = spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_19 = spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_20 = spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_21 = spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_22 = spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_23 = spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_24 = spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_25 = spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_26 = spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_27 = spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_28 = spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_29 = spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_30 = spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_31 = spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_32 = spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_33 = spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_34 = spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_35 = spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_36 = spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_37 = spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_38 = spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_39 = spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_40 = spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_41 = spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_42 = spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_43 = spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_44 = spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_45 = spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_46 = spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_47 = spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_48 = spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_49 = spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_50 = spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_51 = spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_52 = spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_53 = spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_54 = spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_55 = spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_56 = spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_57 = spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_58 = spriteVisibleRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_59 = spriteVisibleRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_60 = spriteVisibleRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_61 = spriteVisibleRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_62 = spriteVisibleRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_63 = spriteVisibleRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_64 = spriteVisibleRegs_64; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_65 = spriteVisibleRegs_65; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_66 = spriteVisibleRegs_66; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_67 = spriteVisibleRegs_67; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_68 = spriteVisibleRegs_68; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_69 = spriteVisibleRegs_69; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_70 = spriteVisibleRegs_70; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_71 = spriteVisibleRegs_71; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_72 = spriteVisibleRegs_72; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_73 = spriteVisibleRegs_73; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_74 = spriteVisibleRegs_74; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_75 = spriteVisibleRegs_75; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_76 = spriteVisibleRegs_76; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_77 = spriteVisibleRegs_77; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_78 = spriteVisibleRegs_78; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_79 = spriteVisibleRegs_79; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_80 = spriteVisibleRegs_80; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_81 = spriteVisibleRegs_81; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_82 = spriteVisibleRegs_82; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_83 = spriteVisibleRegs_83; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_84 = spriteVisibleRegs_84; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_85 = spriteVisibleRegs_85; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_86 = spriteVisibleRegs_86; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_87 = spriteVisibleRegs_87; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_88 = spriteVisibleRegs_88; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_89 = spriteVisibleRegs_89; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_90 = spriteVisibleRegs_90; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_91 = spriteVisibleRegs_91; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_92 = spriteVisibleRegs_92; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_93 = spriteVisibleRegs_93; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_94 = spriteVisibleRegs_94; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_95 = spriteVisibleRegs_95; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_96 = spriteVisibleRegs_96; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_97 = spriteVisibleRegs_97; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_98 = spriteVisibleRegs_98; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteVisible_99 = spriteVisibleRegs_99; // @[\\src\\main\\scala\\GameLogic.scala 185:25]
  assign io_spriteScaleUpHorizontal_16 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1840; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_17 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1845; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_18 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1850; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_19 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1855; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_20 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1860; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_21 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1865; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_22 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1870; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_23 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1875; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_24 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1880; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_25 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1885; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_26 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1840; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_27 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1845; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_28 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1850; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_29 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1855; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_30 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1860; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_31 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1865; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_32 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1870; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_33 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1875; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_34 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1880; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_35 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1885; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_36 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1840; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_37 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1845; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_38 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1850; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_39 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1855; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_40 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1860; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_41 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1865; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_42 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1870; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_43 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1875; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_44 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1880; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_45 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1885; // @[\\src\\main\\scala\\GameLogic.scala 346:20 195:35]
  assign io_spriteScaleUpHorizontal_58 = sprite58ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 201:34]
  assign io_spriteScaleUpHorizontal_59 = sprite59ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 203:34]
  assign io_spriteScaleUpHorizontal_60 = sprite60ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 205:34]
  assign io_spriteScaleUpVertical_16 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1840; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_17 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1845; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_18 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1850; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_19 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1855; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_20 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1860; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_21 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1865; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_22 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1870; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_23 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1875; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_24 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1880; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_25 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1885; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_26 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1840; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_27 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1845; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_28 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1850; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_29 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1855; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_30 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1860; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_31 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1865; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_32 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1870; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_33 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1875; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_34 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1880; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_35 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1885; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_36 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1840; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_37 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1845; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_38 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1850; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_39 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1855; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_40 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1860; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_41 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1865; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_42 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1870; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_43 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1875; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_44 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1880; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_45 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1885; // @[\\src\\main\\scala\\GameLogic.scala 346:20 196:33]
  assign io_spriteScaleUpVertical_58 = sprite58ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 202:32]
  assign io_spriteScaleUpVertical_59 = sprite59ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 204:32]
  assign io_spriteScaleUpVertical_60 = sprite60ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 206:32]
  assign io_viewBoxX = viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 213:15]
  assign io_viewBoxY = viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 214:15]
  assign io_frameUpdateDone = 3'h0 == stateReg ? 1'h0 : _GEN_2100; // @[\\src\\main\\scala\\GameLogic.scala 346:20 100:22]
  assign difficulty_clock = clock;
  assign difficulty_reset = reset;
  assign difficulty_io_level = lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 220:23]
  assign difficulty_io_resetSpeed = gameOverReturnPressed; // @[\\src\\main\\scala\\GameLogic.scala 240:28]
  assign lfsr_clock = clock;
  assign lfsr_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 113:25]
      stateReg <= 3'h0; // @[\\src\\main\\scala\\GameLogic.scala 113:25]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          stateReg <= 3'h2; // @[\\src\\main\\scala\\GameLogic.scala 352:20]
        end else begin
          stateReg <= _GEN_198;
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (livesReg > 3'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 694:28]
        stateReg <= 3'h2; // @[\\src\\main\\scala\\GameLogic.scala 695:18]
      end else begin
        stateReg <= _GEN_1575;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      stateReg <= _GEN_1680;
    end else begin
      stateReg <= _GEN_1781;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_3 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_3 <= _GEN_0;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_3 <= _GEN_0;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_3 <= _GEN_0;
    end else begin
      spriteXRegs_3 <= _GEN_1783;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_7 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_7 <= 11'sh100; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_8 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_8 <= 11'sh100; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_9 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_9 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_10 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_10 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_11 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_11 <= 11'sh160; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_12 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_12 <= 11'sh160; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_13 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_13 <= _GEN_14;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteXRegs_13 <= _GEN_469;
      end else begin
        spriteXRegs_13 <= _GEN_14;
      end
    end else begin
      spriteXRegs_13 <= _GEN_14;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_14 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_14 <= _GEN_16;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_14 <= _GEN_16;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_14 <= _GEN_16;
    end else begin
      spriteXRegs_14 <= _GEN_1766;
    end
    spriteXRegs_16 <= _GEN_2775[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_17 <= _GEN_2777[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_18 <= _GEN_2779[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_19 <= _GEN_2781[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_20 <= _GEN_2783[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_21 <= _GEN_2785[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_22 <= _GEN_2787[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_23 <= _GEN_2789[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_24 <= _GEN_2791[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_25 <= _GEN_2793[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_26 <= _GEN_2795[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_27 <= _GEN_2797[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_28 <= _GEN_2799[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_29 <= _GEN_2801[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_30 <= _GEN_2803[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_31 <= _GEN_2805[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_32 <= _GEN_2807[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_33 <= _GEN_2809[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_34 <= _GEN_2811[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_35 <= _GEN_2813[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_36 <= _GEN_2815[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_37 <= _GEN_2817[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_38 <= _GEN_2819[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_39 <= _GEN_2821[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_40 <= _GEN_2823[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_41 <= _GEN_2825[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_42 <= _GEN_2827[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_43 <= _GEN_2829[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_44 <= _GEN_2831[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_45 <= _GEN_2833[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_46 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_46 <= 11'she0; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_47 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_47 <= 11'sh100; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_48 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_48 <= 11'sh120; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_49 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_49 <= 11'sh140; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_50 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_50 <= 11'sh160; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_51 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_51 <= 11'sh180; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_52 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_52 <= 11'sh110; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_53 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_53 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_54 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_54 <= 11'sh150; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_55 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_55 <= 11'sh110; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_56 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_56 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_57 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_57 <= 11'sh150; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_58 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_58 <= _GEN_102;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 604:29]
        spriteXRegs_58 <= spriteXRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 605:25]
      end else begin
        spriteXRegs_58 <= _GEN_1637;
      end
    end else begin
      spriteXRegs_58 <= _GEN_102;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_59 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_59 <= _GEN_104;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 604:29]
        spriteXRegs_59 <= spriteXRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 607:25]
      end else begin
        spriteXRegs_59 <= _GEN_1638;
      end
    end else begin
      spriteXRegs_59 <= _GEN_104;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_60 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteXRegs_60 <= _GEN_106;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 604:29]
        spriteXRegs_60 <= spriteXRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 609:25]
      end else begin
        spriteXRegs_60 <= _GEN_1639;
      end
    end else begin
      spriteXRegs_60 <= _GEN_106;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_61 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_61 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_62 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_62 <= 11'sh3c; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_63 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_63 <= 11'sh64; // @[\\src\\main\\scala\\GameLogic.scala 169:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_3 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_3 <= _GEN_1;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_3 <= _GEN_1;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_3 <= _GEN_1;
    end else begin
      spriteYRegs_3 <= _GEN_1782;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_7 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_7 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_8 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_8 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_9 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_9 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_10 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_10 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_11 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_11 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_12 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_12 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_13 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_13 <= _GEN_15;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_13 <= _GEN_467;
      end else begin
        spriteYRegs_13 <= _GEN_15;
      end
    end else begin
      spriteYRegs_13 <= _GEN_15;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_14 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_14 <= _GEN_17;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_14 <= _GEN_17;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_14 <= _GEN_17;
    end else begin
      spriteYRegs_14 <= _GEN_1767;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_16 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_16 <= _GEN_19;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_16 <= _GEN_317;
      end else begin
        spriteYRegs_16 <= _GEN_19;
      end
    end else begin
      spriteYRegs_16 <= _GEN_19;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_17 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_17 <= _GEN_21;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_17 <= _GEN_322;
      end else begin
        spriteYRegs_17 <= _GEN_21;
      end
    end else begin
      spriteYRegs_17 <= _GEN_21;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_18 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_18 <= _GEN_23;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_18 <= _GEN_327;
      end else begin
        spriteYRegs_18 <= _GEN_23;
      end
    end else begin
      spriteYRegs_18 <= _GEN_23;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_19 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_19 <= _GEN_25;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_19 <= _GEN_332;
      end else begin
        spriteYRegs_19 <= _GEN_25;
      end
    end else begin
      spriteYRegs_19 <= _GEN_25;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_20 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_20 <= _GEN_27;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_20 <= _GEN_337;
      end else begin
        spriteYRegs_20 <= _GEN_27;
      end
    end else begin
      spriteYRegs_20 <= _GEN_27;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_21 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_21 <= _GEN_29;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_21 <= _GEN_342;
      end else begin
        spriteYRegs_21 <= _GEN_29;
      end
    end else begin
      spriteYRegs_21 <= _GEN_29;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_22 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_22 <= _GEN_31;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_22 <= _GEN_347;
      end else begin
        spriteYRegs_22 <= _GEN_31;
      end
    end else begin
      spriteYRegs_22 <= _GEN_31;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_23 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_23 <= _GEN_33;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_23 <= _GEN_352;
      end else begin
        spriteYRegs_23 <= _GEN_33;
      end
    end else begin
      spriteYRegs_23 <= _GEN_33;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_24 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_24 <= _GEN_35;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_24 <= _GEN_357;
      end else begin
        spriteYRegs_24 <= _GEN_35;
      end
    end else begin
      spriteYRegs_24 <= _GEN_35;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_25 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_25 <= _GEN_37;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_25 <= _GEN_362;
      end else begin
        spriteYRegs_25 <= _GEN_37;
      end
    end else begin
      spriteYRegs_25 <= _GEN_37;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_26 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_26 <= _GEN_39;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_26 <= _GEN_367;
      end else begin
        spriteYRegs_26 <= _GEN_39;
      end
    end else begin
      spriteYRegs_26 <= _GEN_39;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_27 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_27 <= _GEN_41;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_27 <= _GEN_372;
      end else begin
        spriteYRegs_27 <= _GEN_41;
      end
    end else begin
      spriteYRegs_27 <= _GEN_41;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_28 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_28 <= _GEN_43;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_28 <= _GEN_377;
      end else begin
        spriteYRegs_28 <= _GEN_43;
      end
    end else begin
      spriteYRegs_28 <= _GEN_43;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_29 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_29 <= _GEN_45;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_29 <= _GEN_382;
      end else begin
        spriteYRegs_29 <= _GEN_45;
      end
    end else begin
      spriteYRegs_29 <= _GEN_45;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_30 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_30 <= _GEN_47;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_30 <= _GEN_387;
      end else begin
        spriteYRegs_30 <= _GEN_47;
      end
    end else begin
      spriteYRegs_30 <= _GEN_47;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_31 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_31 <= _GEN_49;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_31 <= _GEN_392;
      end else begin
        spriteYRegs_31 <= _GEN_49;
      end
    end else begin
      spriteYRegs_31 <= _GEN_49;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_32 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_32 <= _GEN_51;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_32 <= _GEN_397;
      end else begin
        spriteYRegs_32 <= _GEN_51;
      end
    end else begin
      spriteYRegs_32 <= _GEN_51;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_33 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_33 <= _GEN_53;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_33 <= _GEN_402;
      end else begin
        spriteYRegs_33 <= _GEN_53;
      end
    end else begin
      spriteYRegs_33 <= _GEN_53;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_34 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_34 <= _GEN_55;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_34 <= _GEN_407;
      end else begin
        spriteYRegs_34 <= _GEN_55;
      end
    end else begin
      spriteYRegs_34 <= _GEN_55;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_35 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_35 <= _GEN_57;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_35 <= _GEN_412;
      end else begin
        spriteYRegs_35 <= _GEN_57;
      end
    end else begin
      spriteYRegs_35 <= _GEN_57;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_36 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_36 <= _GEN_59;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_36 <= _GEN_417;
      end else begin
        spriteYRegs_36 <= _GEN_59;
      end
    end else begin
      spriteYRegs_36 <= _GEN_59;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_37 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_37 <= _GEN_61;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_37 <= _GEN_422;
      end else begin
        spriteYRegs_37 <= _GEN_61;
      end
    end else begin
      spriteYRegs_37 <= _GEN_61;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_38 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_38 <= _GEN_63;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_38 <= _GEN_427;
      end else begin
        spriteYRegs_38 <= _GEN_63;
      end
    end else begin
      spriteYRegs_38 <= _GEN_63;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_39 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_39 <= _GEN_65;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_39 <= _GEN_432;
      end else begin
        spriteYRegs_39 <= _GEN_65;
      end
    end else begin
      spriteYRegs_39 <= _GEN_65;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_40 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_40 <= _GEN_67;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_40 <= _GEN_437;
      end else begin
        spriteYRegs_40 <= _GEN_67;
      end
    end else begin
      spriteYRegs_40 <= _GEN_67;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_41 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_41 <= _GEN_69;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_41 <= _GEN_442;
      end else begin
        spriteYRegs_41 <= _GEN_69;
      end
    end else begin
      spriteYRegs_41 <= _GEN_69;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_42 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_42 <= _GEN_71;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_42 <= _GEN_447;
      end else begin
        spriteYRegs_42 <= _GEN_71;
      end
    end else begin
      spriteYRegs_42 <= _GEN_71;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_43 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_43 <= _GEN_73;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_43 <= _GEN_452;
      end else begin
        spriteYRegs_43 <= _GEN_73;
      end
    end else begin
      spriteYRegs_43 <= _GEN_73;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_44 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_44 <= _GEN_75;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_44 <= _GEN_457;
      end else begin
        spriteYRegs_44 <= _GEN_75;
      end
    end else begin
      spriteYRegs_44 <= _GEN_75;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_45 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_45 <= _GEN_77;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        spriteYRegs_45 <= _GEN_462;
      end else begin
        spriteYRegs_45 <= _GEN_77;
      end
    end else begin
      spriteYRegs_45 <= _GEN_77;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_46 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_46 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_47 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_47 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_48 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_48 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_49 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_49 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_50 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_50 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_51 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_51 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_52 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_52 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_53 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_53 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_54 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_54 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_55 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_55 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_56 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_56 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_57 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_57 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_58 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_58 <= _GEN_103;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 604:29]
        spriteYRegs_58 <= spriteYRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 606:25]
      end else begin
        spriteYRegs_58 <= _GEN_1640;
      end
    end else begin
      spriteYRegs_58 <= _GEN_103;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_59 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_59 <= _GEN_105;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 604:29]
        spriteYRegs_59 <= spriteYRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 608:25]
      end else begin
        spriteYRegs_59 <= _GEN_1641;
      end
    end else begin
      spriteYRegs_59 <= _GEN_105;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_60 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteYRegs_60 <= _GEN_107;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 604:29]
        spriteYRegs_60 <= spriteYRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 610:25]
      end else begin
        spriteYRegs_60 <= _GEN_1642;
      end
    end else begin
      spriteYRegs_60 <= _GEN_107;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_61 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_61 <= 10'sh14; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_62 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_62 <= 10'sh14; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_63 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_63 <= 10'sh14; // @[\\src\\main\\scala\\GameLogic.scala 170:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_3 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        spriteVisibleRegs_3 <= _GEN_211;
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_3 <= _GEN_709;
      end else begin
        spriteVisibleRegs_3 <= _GEN_1319;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_3 <= _GEN_1681;
    end else begin
      spriteVisibleRegs_3 <= _GEN_1768;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_4 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_4 <= _GEN_710;
        end else begin
          spriteVisibleRegs_4 <= _GEN_1320;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_5 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_5 <= _GEN_711;
        end else begin
          spriteVisibleRegs_5 <= _GEN_1321;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_6 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_6 <= _GEN_712;
        end else begin
          spriteVisibleRegs_6 <= _GEN_1322;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_7 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_7 <= _GEN_713;
        end else begin
          spriteVisibleRegs_7 <= _GEN_1323;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        spriteVisibleRegs_7 <= _GEN_1682;
      end else begin
        spriteVisibleRegs_7 <= _GEN_1769;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_8 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_8 <= _GEN_714;
        end else begin
          spriteVisibleRegs_8 <= _GEN_1324;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        spriteVisibleRegs_8 <= _GEN_1683;
      end else begin
        spriteVisibleRegs_8 <= _GEN_1770;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_9 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_9 <= _GEN_715;
        end else begin
          spriteVisibleRegs_9 <= _GEN_1325;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        spriteVisibleRegs_9 <= _GEN_1684;
      end else begin
        spriteVisibleRegs_9 <= _GEN_1771;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_10 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_10 <= _GEN_716;
        end else begin
          spriteVisibleRegs_10 <= _GEN_1326;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        spriteVisibleRegs_10 <= _GEN_1685;
      end else begin
        spriteVisibleRegs_10 <= _GEN_1772;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_11 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_11 <= _GEN_717;
        end else begin
          spriteVisibleRegs_11 <= _GEN_1327;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        spriteVisibleRegs_11 <= _GEN_1686;
      end else begin
        spriteVisibleRegs_11 <= _GEN_1773;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_12 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_12 <= _GEN_718;
        end else begin
          spriteVisibleRegs_12 <= _GEN_1328;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        spriteVisibleRegs_12 <= _GEN_1687;
      end else begin
        spriteVisibleRegs_12 <= _GEN_1774;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_13 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T_792) begin // @[\\src\\main\\scala\\GameLogic.scala 550:9]
          spriteVisibleRegs_13 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 551:31]
        end else begin
          spriteVisibleRegs_13 <= _GEN_1431;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_14 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_14 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:27]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 565:24]
        spriteVisibleRegs_14 <= _GEN_1566;
      end else begin
        spriteVisibleRegs_14 <= _GEN_1432;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_14 <= _GEN_1775;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_15 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_15 <= _GEN_721;
        end else begin
          spriteVisibleRegs_15 <= _GEN_1331;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_16 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_16 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_16 <= _GEN_722;
      end else begin
        spriteVisibleRegs_16 <= _GEN_1332;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_17 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_17 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_17 <= _GEN_723;
      end else begin
        spriteVisibleRegs_17 <= _GEN_1333;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_18 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_18 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_18 <= _GEN_724;
      end else begin
        spriteVisibleRegs_18 <= _GEN_1334;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_19 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_19 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_19 <= _GEN_725;
      end else begin
        spriteVisibleRegs_19 <= _GEN_1335;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_20 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_20 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_20 <= _GEN_726;
      end else begin
        spriteVisibleRegs_20 <= _GEN_1336;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_21 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_21 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_21 <= _GEN_727;
      end else begin
        spriteVisibleRegs_21 <= _GEN_1337;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_22 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_22 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_22 <= _GEN_728;
      end else begin
        spriteVisibleRegs_22 <= _GEN_1338;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_23 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_23 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_23 <= _GEN_729;
      end else begin
        spriteVisibleRegs_23 <= _GEN_1339;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_24 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_24 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_24 <= _GEN_730;
      end else begin
        spriteVisibleRegs_24 <= _GEN_1340;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_25 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_25 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_25 <= _GEN_731;
      end else begin
        spriteVisibleRegs_25 <= _GEN_1341;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_26 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_26 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_26 <= _GEN_732;
      end else begin
        spriteVisibleRegs_26 <= _GEN_1342;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_27 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_27 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_27 <= _GEN_733;
      end else begin
        spriteVisibleRegs_27 <= _GEN_1343;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_28 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_28 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_28 <= _GEN_734;
      end else begin
        spriteVisibleRegs_28 <= _GEN_1344;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_29 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_29 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_29 <= _GEN_735;
      end else begin
        spriteVisibleRegs_29 <= _GEN_1345;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_30 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_30 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_30 <= _GEN_736;
      end else begin
        spriteVisibleRegs_30 <= _GEN_1346;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_31 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_31 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_31 <= _GEN_737;
      end else begin
        spriteVisibleRegs_31 <= _GEN_1347;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_32 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_32 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_32 <= _GEN_738;
      end else begin
        spriteVisibleRegs_32 <= _GEN_1348;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_33 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_33 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_33 <= _GEN_739;
      end else begin
        spriteVisibleRegs_33 <= _GEN_1349;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_34 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_34 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_34 <= _GEN_740;
      end else begin
        spriteVisibleRegs_34 <= _GEN_1350;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_35 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_35 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_35 <= _GEN_741;
      end else begin
        spriteVisibleRegs_35 <= _GEN_1351;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_36 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_36 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_36 <= _GEN_742;
      end else begin
        spriteVisibleRegs_36 <= _GEN_1352;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_37 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_37 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_37 <= _GEN_743;
      end else begin
        spriteVisibleRegs_37 <= _GEN_1353;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_38 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_38 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_38 <= _GEN_744;
      end else begin
        spriteVisibleRegs_38 <= _GEN_1354;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_39 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_39 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_39 <= _GEN_745;
      end else begin
        spriteVisibleRegs_39 <= _GEN_1355;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_40 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_40 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_40 <= _GEN_746;
      end else begin
        spriteVisibleRegs_40 <= _GEN_1356;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_41 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_41 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_41 <= _GEN_747;
      end else begin
        spriteVisibleRegs_41 <= _GEN_1357;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_42 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_42 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_42 <= _GEN_748;
      end else begin
        spriteVisibleRegs_42 <= _GEN_1358;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_43 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_43 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_43 <= _GEN_749;
      end else begin
        spriteVisibleRegs_43 <= _GEN_1359;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_44 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_44 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_44 <= _GEN_750;
      end else begin
        spriteVisibleRegs_44 <= _GEN_1360;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_45 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_45 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 310:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_45 <= _GEN_751;
      end else begin
        spriteVisibleRegs_45 <= _GEN_1361;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_46 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_46 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_46 <= _GEN_752;
      end else begin
        spriteVisibleRegs_46 <= _GEN_1362;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_46 <= _GEN_1784;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_47 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_47 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_47 <= _GEN_753;
      end else begin
        spriteVisibleRegs_47 <= _GEN_1363;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_47 <= _GEN_1785;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_48 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_48 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_48 <= _GEN_754;
      end else begin
        spriteVisibleRegs_48 <= _GEN_1364;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_48 <= _GEN_1786;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_49 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_49 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_49 <= _GEN_755;
      end else begin
        spriteVisibleRegs_49 <= _GEN_1365;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_49 <= _GEN_1787;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_50 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_50 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_50 <= _GEN_756;
      end else begin
        spriteVisibleRegs_50 <= _GEN_1366;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_50 <= _GEN_1788;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_51 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_51 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_51 <= _GEN_757;
      end else begin
        spriteVisibleRegs_51 <= _GEN_1367;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_51 <= _GEN_1789;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_52 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_52 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_52 <= _GEN_758;
      end else begin
        spriteVisibleRegs_52 <= _GEN_1368;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_52 <= _GEN_1790;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_53 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_53 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_53 <= _GEN_759;
      end else begin
        spriteVisibleRegs_53 <= _GEN_1369;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_53 <= _GEN_1791;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_54 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_54 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_54 <= _GEN_760;
      end else begin
        spriteVisibleRegs_54 <= _GEN_1370;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_54 <= _GEN_1792;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_55 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_55 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_55 <= _GEN_761;
      end else begin
        spriteVisibleRegs_55 <= _GEN_1371;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_55 <= _GEN_1793;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_56 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_56 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_56 <= _GEN_762;
      end else begin
        spriteVisibleRegs_56 <= _GEN_1372;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_56 <= _GEN_1794;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_57 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spriteVisibleRegs_57 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 315:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_57 <= _GEN_763;
      end else begin
        spriteVisibleRegs_57 <= _GEN_1373;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_57 <= _GEN_1795;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_58 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        spriteVisibleRegs_58 <= _T_83;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_59 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        spriteVisibleRegs_59 <= _T_83;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_60 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        spriteVisibleRegs_60 <= _T_83;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_61 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_61 <= _GEN_195;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_61 <= _GEN_767;
      end else begin
        spriteVisibleRegs_61 <= _GEN_1377;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_61 <= _GEN_195;
    end else begin
      spriteVisibleRegs_61 <= _GEN_1776;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_62 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_62 <= _GEN_196;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_62 <= _GEN_768;
      end else begin
        spriteVisibleRegs_62 <= _GEN_1378;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_62 <= _GEN_196;
    end else begin
      spriteVisibleRegs_62 <= _GEN_1777;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_63 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_63 <= _GEN_197;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spriteVisibleRegs_63 <= _GEN_769;
      end else begin
        spriteVisibleRegs_63 <= _GEN_1379;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spriteVisibleRegs_63 <= _GEN_197;
    end else begin
      spriteVisibleRegs_63 <= _GEN_1778;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_64 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_64 <= _GEN_770;
        end else begin
          spriteVisibleRegs_64 <= _GEN_1380;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_65 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_65 <= _GEN_771;
        end else begin
          spriteVisibleRegs_65 <= _GEN_1381;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_66 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_66 <= _GEN_772;
        end else begin
          spriteVisibleRegs_66 <= _GEN_1382;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_67 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_67 <= _GEN_773;
        end else begin
          spriteVisibleRegs_67 <= _GEN_1383;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_68 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_68 <= _GEN_774;
        end else begin
          spriteVisibleRegs_68 <= _GEN_1384;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_69 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_69 <= _GEN_775;
        end else begin
          spriteVisibleRegs_69 <= _GEN_1385;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_70 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_70 <= _GEN_776;
        end else begin
          spriteVisibleRegs_70 <= _GEN_1386;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_71 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_71 <= _GEN_777;
        end else begin
          spriteVisibleRegs_71 <= _GEN_1387;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_72 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_72 <= _GEN_778;
        end else begin
          spriteVisibleRegs_72 <= _GEN_1388;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_73 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_73 <= _GEN_779;
        end else begin
          spriteVisibleRegs_73 <= _GEN_1389;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_74 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_74 <= _GEN_780;
        end else begin
          spriteVisibleRegs_74 <= _GEN_1390;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_75 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_75 <= _GEN_781;
        end else begin
          spriteVisibleRegs_75 <= _GEN_1391;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_76 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_76 <= _GEN_782;
        end else begin
          spriteVisibleRegs_76 <= _GEN_1392;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_77 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_77 <= _GEN_783;
        end else begin
          spriteVisibleRegs_77 <= _GEN_1393;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_78 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_78 <= _GEN_784;
        end else begin
          spriteVisibleRegs_78 <= _GEN_1394;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_79 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_79 <= _GEN_785;
        end else begin
          spriteVisibleRegs_79 <= _GEN_1395;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_80 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_80 <= _GEN_786;
        end else begin
          spriteVisibleRegs_80 <= _GEN_1396;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_81 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_81 <= _GEN_787;
        end else begin
          spriteVisibleRegs_81 <= _GEN_1397;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_82 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_82 <= _GEN_788;
        end else begin
          spriteVisibleRegs_82 <= _GEN_1398;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_83 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_83 <= _GEN_789;
        end else begin
          spriteVisibleRegs_83 <= _GEN_1399;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_84 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_84 <= _GEN_790;
        end else begin
          spriteVisibleRegs_84 <= _GEN_1400;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_85 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_85 <= _GEN_791;
        end else begin
          spriteVisibleRegs_85 <= _GEN_1401;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_86 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_86 <= _GEN_792;
        end else begin
          spriteVisibleRegs_86 <= _GEN_1402;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_87 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_87 <= _GEN_793;
        end else begin
          spriteVisibleRegs_87 <= _GEN_1403;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_88 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_88 <= _GEN_794;
        end else begin
          spriteVisibleRegs_88 <= _GEN_1404;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_89 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_89 <= _GEN_795;
        end else begin
          spriteVisibleRegs_89 <= _GEN_1405;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_90 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_90 <= _GEN_796;
        end else begin
          spriteVisibleRegs_90 <= _GEN_1406;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_91 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_91 <= _GEN_797;
        end else begin
          spriteVisibleRegs_91 <= _GEN_1407;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_92 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_92 <= _GEN_798;
        end else begin
          spriteVisibleRegs_92 <= _GEN_1408;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_93 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_93 <= _GEN_799;
        end else begin
          spriteVisibleRegs_93 <= _GEN_1409;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_94 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_94 <= _GEN_800;
        end else begin
          spriteVisibleRegs_94 <= _GEN_1410;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_95 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_95 <= _GEN_801;
        end else begin
          spriteVisibleRegs_95 <= _GEN_1411;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_96 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_96 <= _GEN_802;
        end else begin
          spriteVisibleRegs_96 <= _GEN_1412;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_97 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_97 <= _GEN_803;
        end else begin
          spriteVisibleRegs_97 <= _GEN_1413;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_98 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_98 <= _GEN_804;
        end else begin
          spriteVisibleRegs_98 <= _GEN_1414;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_99 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
          spriteVisibleRegs_99 <= _GEN_805;
        end else begin
          spriteVisibleRegs_99 <= _GEN_1415;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_0 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_0 <= _GEN_418;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_1 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_1 <= _GEN_423;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_2 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_2 <= _GEN_428;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_3 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_3 <= _GEN_433;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_4 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_4 <= _GEN_438;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_5 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_5 <= _GEN_443;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_6 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_6 <= _GEN_448;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_7 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_7 <= _GEN_453;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_8 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_8 <= _GEN_458;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_9 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
          spriteScaleTypeRegs_9 <= _GEN_463;
        end
      end
    end
    initializePositions <= reset | _GEN_2112; // @[\\src\\main\\scala\\GameLogic.scala 130:{36,36}]
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 176:42]
      sprite58ScaleUpHorizontal <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 176:42]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        sprite58ScaleUpHorizontal <= _GEN_1650;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 177:40]
      sprite58ScaleUpVertical <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 177:40]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        sprite58ScaleUpVertical <= _GEN_1653;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 178:42]
      sprite59ScaleUpHorizontal <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 178:42]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        sprite59ScaleUpHorizontal <= _GEN_1651;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 179:40]
      sprite59ScaleUpVertical <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 179:40]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        sprite59ScaleUpVertical <= _GEN_1654;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 180:42]
      sprite60ScaleUpHorizontal <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 180:42]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        sprite60ScaleUpHorizontal <= _GEN_1652;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 181:40]
      sprite60ScaleUpVertical <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 181:40]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        sprite60ScaleUpVertical <= _GEN_1655;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 209:28]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 209:28]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
          viewBoxXReg <= _GEN_1779;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 210:28]
      viewBoxYReg <= 9'h0; // @[\\src\\main\\scala\\GameLogic.scala 210:28]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
          viewBoxYReg <= _GEN_1780;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 219:23]
      lvlReg <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 219:23]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          lvlReg <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 291:12]
        end
      end
    end else if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        lvlReg <= _GEN_1688;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 231:25]
      livesReg <= 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 231:25]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          livesReg <= 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 292:14]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 565:24]
        livesReg <= _GEN_1567;
      end else begin
        livesReg <= _GEN_1555;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 234:29]
      extraLifeCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 234:29]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          extraLifeCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 296:18]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 369:29]
        extraLifeCnt <= _GEN_468;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 237:38]
      gameOverReturnPressed <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 237:38]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          gameOverReturnPressed <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 351:33]
        end
      end
    end else if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
        gameOverReturnPressed <= _GEN_1796;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 243:34]
      spawnDelayCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 243:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          spawnDelayCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 294:23]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        spawnDelayCounter <= _GEN_807;
      end else begin
        spawnDelayCounter <= _GEN_1417;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      spawnDelayCounter <= _GEN_1765;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 244:34]
      nextSpriteToSpawn <= 6'h0; // @[\\src\\main\\scala\\GameLogic.scala 244:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          nextSpriteToSpawn <= 6'h0; // @[\\src\\main\\scala\\GameLogic.scala 295:23]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 460:28]
        nextSpriteToSpawn <= _GEN_806;
      end else begin
        nextSpriteToSpawn <= _GEN_1416;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      nextSpriteToSpawn <= _GEN_1764;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 247:24]
      starCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 247:24]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          starCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 297:13]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 604:29]
        starCnt <= _starCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 617:17]
      end else begin
        starCnt <= _GEN_1643;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 250:34]
      collisionDetected <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 250:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          collisionDetected <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 298:23]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 565:24]
        collisionDetected <= _GEN_1569;
      end else begin
        collisionDetected <= _GEN_1552;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 251:29]
      blinkCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 251:29]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          blinkCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 300:18]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 565:24]
        blinkCounter <= _GEN_1561;
      end else begin
        blinkCounter <= _GEN_1557;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 252:27]
      blinkTimes <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 252:27]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          blinkTimes <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:16]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 565:24]
        blinkTimes <= _GEN_1562;
      end else begin
        blinkTimes <= _GEN_1558;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 253:27]
      isBlinking <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 253:27]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 348:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 349:37]
          isBlinking <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 299:16]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 346:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 565:24]
        isBlinking <= _GEN_1565;
      end else begin
        isBlinking <= _GEN_1556;
      end
    end
    spriteXRegs_58_REG <= $signed(spriteXRegs_59) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 605:52]
    spriteYRegs_58_REG <= $signed(spriteYRegs_59) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 606:52]
    spriteXRegs_59_REG <= $signed(spriteXRegs_60) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 607:52]
    spriteYRegs_59_REG <= $signed(spriteYRegs_60) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 608:52]
    spriteXRegs_60_REG <= $signed(spriteXRegs_58) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 609:52]
    spriteYRegs_60_REG <= $signed(spriteYRegs_58) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 610:52]
    spriteXRegs_58_REG_1 <= $signed(spriteXRegs_59) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 633:52]
    spriteYRegs_58_REG_1 <= $signed(spriteYRegs_59) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 634:52]
    spriteXRegs_59_REG_1 <= $signed(spriteXRegs_60) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 635:52]
    spriteYRegs_59_REG_1 <= $signed(spriteYRegs_60) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 636:52]
    spriteXRegs_60_REG_1 <= $signed(spriteXRegs_58) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 637:52]
    spriteYRegs_60_REG_1 <= $signed(spriteYRegs_58) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 638:52]
    spriteXRegs_58_REG_2 <= $signed(spriteXRegs_59) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 661:52]
    spriteYRegs_58_REG_2 <= $signed(spriteYRegs_59) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 662:52]
    spriteXRegs_59_REG_2 <= $signed(spriteXRegs_60) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 663:52]
    spriteYRegs_59_REG_2 <= $signed(spriteYRegs_60) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 664:52]
    spriteXRegs_60_REG_2 <= $signed(spriteXRegs_58) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 665:52]
    spriteYRegs_60_REG_2 <= $signed(spriteYRegs_58) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 666:52]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  spriteXRegs_3 = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  spriteXRegs_7 = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  spriteXRegs_8 = _RAND_3[10:0];
  _RAND_4 = {1{`RANDOM}};
  spriteXRegs_9 = _RAND_4[10:0];
  _RAND_5 = {1{`RANDOM}};
  spriteXRegs_10 = _RAND_5[10:0];
  _RAND_6 = {1{`RANDOM}};
  spriteXRegs_11 = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  spriteXRegs_12 = _RAND_7[10:0];
  _RAND_8 = {1{`RANDOM}};
  spriteXRegs_13 = _RAND_8[10:0];
  _RAND_9 = {1{`RANDOM}};
  spriteXRegs_14 = _RAND_9[10:0];
  _RAND_10 = {1{`RANDOM}};
  spriteXRegs_16 = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  spriteXRegs_17 = _RAND_11[10:0];
  _RAND_12 = {1{`RANDOM}};
  spriteXRegs_18 = _RAND_12[10:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXRegs_19 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXRegs_20 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXRegs_21 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXRegs_22 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXRegs_23 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXRegs_24 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXRegs_25 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteXRegs_26 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  spriteXRegs_27 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  spriteXRegs_28 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  spriteXRegs_29 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  spriteXRegs_30 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  spriteXRegs_31 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  spriteXRegs_32 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  spriteXRegs_33 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  spriteXRegs_34 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  spriteXRegs_35 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  spriteXRegs_36 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  spriteXRegs_37 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  spriteXRegs_38 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  spriteXRegs_39 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  spriteXRegs_40 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  spriteXRegs_41 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  spriteXRegs_42 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  spriteXRegs_43 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  spriteXRegs_44 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  spriteXRegs_45 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  spriteXRegs_46 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  spriteXRegs_47 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  spriteXRegs_48 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  spriteXRegs_49 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  spriteXRegs_50 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  spriteXRegs_51 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  spriteXRegs_52 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  spriteXRegs_53 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  spriteXRegs_54 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  spriteXRegs_55 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  spriteXRegs_56 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  spriteXRegs_57 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  spriteXRegs_58 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  spriteXRegs_59 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  spriteXRegs_60 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  spriteXRegs_61 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  spriteXRegs_62 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  spriteXRegs_63 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  spriteYRegs_3 = _RAND_58[9:0];
  _RAND_59 = {1{`RANDOM}};
  spriteYRegs_7 = _RAND_59[9:0];
  _RAND_60 = {1{`RANDOM}};
  spriteYRegs_8 = _RAND_60[9:0];
  _RAND_61 = {1{`RANDOM}};
  spriteYRegs_9 = _RAND_61[9:0];
  _RAND_62 = {1{`RANDOM}};
  spriteYRegs_10 = _RAND_62[9:0];
  _RAND_63 = {1{`RANDOM}};
  spriteYRegs_11 = _RAND_63[9:0];
  _RAND_64 = {1{`RANDOM}};
  spriteYRegs_12 = _RAND_64[9:0];
  _RAND_65 = {1{`RANDOM}};
  spriteYRegs_13 = _RAND_65[9:0];
  _RAND_66 = {1{`RANDOM}};
  spriteYRegs_14 = _RAND_66[9:0];
  _RAND_67 = {1{`RANDOM}};
  spriteYRegs_16 = _RAND_67[9:0];
  _RAND_68 = {1{`RANDOM}};
  spriteYRegs_17 = _RAND_68[9:0];
  _RAND_69 = {1{`RANDOM}};
  spriteYRegs_18 = _RAND_69[9:0];
  _RAND_70 = {1{`RANDOM}};
  spriteYRegs_19 = _RAND_70[9:0];
  _RAND_71 = {1{`RANDOM}};
  spriteYRegs_20 = _RAND_71[9:0];
  _RAND_72 = {1{`RANDOM}};
  spriteYRegs_21 = _RAND_72[9:0];
  _RAND_73 = {1{`RANDOM}};
  spriteYRegs_22 = _RAND_73[9:0];
  _RAND_74 = {1{`RANDOM}};
  spriteYRegs_23 = _RAND_74[9:0];
  _RAND_75 = {1{`RANDOM}};
  spriteYRegs_24 = _RAND_75[9:0];
  _RAND_76 = {1{`RANDOM}};
  spriteYRegs_25 = _RAND_76[9:0];
  _RAND_77 = {1{`RANDOM}};
  spriteYRegs_26 = _RAND_77[9:0];
  _RAND_78 = {1{`RANDOM}};
  spriteYRegs_27 = _RAND_78[9:0];
  _RAND_79 = {1{`RANDOM}};
  spriteYRegs_28 = _RAND_79[9:0];
  _RAND_80 = {1{`RANDOM}};
  spriteYRegs_29 = _RAND_80[9:0];
  _RAND_81 = {1{`RANDOM}};
  spriteYRegs_30 = _RAND_81[9:0];
  _RAND_82 = {1{`RANDOM}};
  spriteYRegs_31 = _RAND_82[9:0];
  _RAND_83 = {1{`RANDOM}};
  spriteYRegs_32 = _RAND_83[9:0];
  _RAND_84 = {1{`RANDOM}};
  spriteYRegs_33 = _RAND_84[9:0];
  _RAND_85 = {1{`RANDOM}};
  spriteYRegs_34 = _RAND_85[9:0];
  _RAND_86 = {1{`RANDOM}};
  spriteYRegs_35 = _RAND_86[9:0];
  _RAND_87 = {1{`RANDOM}};
  spriteYRegs_36 = _RAND_87[9:0];
  _RAND_88 = {1{`RANDOM}};
  spriteYRegs_37 = _RAND_88[9:0];
  _RAND_89 = {1{`RANDOM}};
  spriteYRegs_38 = _RAND_89[9:0];
  _RAND_90 = {1{`RANDOM}};
  spriteYRegs_39 = _RAND_90[9:0];
  _RAND_91 = {1{`RANDOM}};
  spriteYRegs_40 = _RAND_91[9:0];
  _RAND_92 = {1{`RANDOM}};
  spriteYRegs_41 = _RAND_92[9:0];
  _RAND_93 = {1{`RANDOM}};
  spriteYRegs_42 = _RAND_93[9:0];
  _RAND_94 = {1{`RANDOM}};
  spriteYRegs_43 = _RAND_94[9:0];
  _RAND_95 = {1{`RANDOM}};
  spriteYRegs_44 = _RAND_95[9:0];
  _RAND_96 = {1{`RANDOM}};
  spriteYRegs_45 = _RAND_96[9:0];
  _RAND_97 = {1{`RANDOM}};
  spriteYRegs_46 = _RAND_97[9:0];
  _RAND_98 = {1{`RANDOM}};
  spriteYRegs_47 = _RAND_98[9:0];
  _RAND_99 = {1{`RANDOM}};
  spriteYRegs_48 = _RAND_99[9:0];
  _RAND_100 = {1{`RANDOM}};
  spriteYRegs_49 = _RAND_100[9:0];
  _RAND_101 = {1{`RANDOM}};
  spriteYRegs_50 = _RAND_101[9:0];
  _RAND_102 = {1{`RANDOM}};
  spriteYRegs_51 = _RAND_102[9:0];
  _RAND_103 = {1{`RANDOM}};
  spriteYRegs_52 = _RAND_103[9:0];
  _RAND_104 = {1{`RANDOM}};
  spriteYRegs_53 = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  spriteYRegs_54 = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  spriteYRegs_55 = _RAND_106[9:0];
  _RAND_107 = {1{`RANDOM}};
  spriteYRegs_56 = _RAND_107[9:0];
  _RAND_108 = {1{`RANDOM}};
  spriteYRegs_57 = _RAND_108[9:0];
  _RAND_109 = {1{`RANDOM}};
  spriteYRegs_58 = _RAND_109[9:0];
  _RAND_110 = {1{`RANDOM}};
  spriteYRegs_59 = _RAND_110[9:0];
  _RAND_111 = {1{`RANDOM}};
  spriteYRegs_60 = _RAND_111[9:0];
  _RAND_112 = {1{`RANDOM}};
  spriteYRegs_61 = _RAND_112[9:0];
  _RAND_113 = {1{`RANDOM}};
  spriteYRegs_62 = _RAND_113[9:0];
  _RAND_114 = {1{`RANDOM}};
  spriteYRegs_63 = _RAND_114[9:0];
  _RAND_115 = {1{`RANDOM}};
  spriteVisibleRegs_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  spriteVisibleRegs_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  spriteVisibleRegs_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  spriteVisibleRegs_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  spriteVisibleRegs_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  spriteVisibleRegs_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  spriteVisibleRegs_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  spriteVisibleRegs_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  spriteVisibleRegs_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  spriteVisibleRegs_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  spriteVisibleRegs_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  spriteVisibleRegs_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  spriteVisibleRegs_15 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  spriteVisibleRegs_16 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  spriteVisibleRegs_17 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  spriteVisibleRegs_18 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  spriteVisibleRegs_19 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  spriteVisibleRegs_20 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  spriteVisibleRegs_21 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  spriteVisibleRegs_22 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  spriteVisibleRegs_23 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  spriteVisibleRegs_24 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  spriteVisibleRegs_25 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  spriteVisibleRegs_26 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  spriteVisibleRegs_27 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  spriteVisibleRegs_28 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  spriteVisibleRegs_29 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  spriteVisibleRegs_30 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  spriteVisibleRegs_31 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  spriteVisibleRegs_32 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  spriteVisibleRegs_33 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  spriteVisibleRegs_34 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  spriteVisibleRegs_35 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  spriteVisibleRegs_36 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  spriteVisibleRegs_37 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  spriteVisibleRegs_38 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  spriteVisibleRegs_39 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  spriteVisibleRegs_40 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  spriteVisibleRegs_41 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  spriteVisibleRegs_42 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  spriteVisibleRegs_43 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  spriteVisibleRegs_44 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  spriteVisibleRegs_45 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  spriteVisibleRegs_46 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  spriteVisibleRegs_47 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  spriteVisibleRegs_48 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  spriteVisibleRegs_49 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  spriteVisibleRegs_50 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  spriteVisibleRegs_51 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  spriteVisibleRegs_52 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  spriteVisibleRegs_53 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  spriteVisibleRegs_54 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  spriteVisibleRegs_55 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  spriteVisibleRegs_56 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  spriteVisibleRegs_57 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  spriteVisibleRegs_58 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  spriteVisibleRegs_59 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  spriteVisibleRegs_60 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  spriteVisibleRegs_61 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  spriteVisibleRegs_62 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  spriteVisibleRegs_63 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  spriteVisibleRegs_64 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  spriteVisibleRegs_65 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  spriteVisibleRegs_66 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  spriteVisibleRegs_67 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  spriteVisibleRegs_68 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  spriteVisibleRegs_69 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  spriteVisibleRegs_70 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  spriteVisibleRegs_71 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  spriteVisibleRegs_72 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  spriteVisibleRegs_73 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  spriteVisibleRegs_74 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  spriteVisibleRegs_75 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  spriteVisibleRegs_76 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  spriteVisibleRegs_77 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  spriteVisibleRegs_78 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  spriteVisibleRegs_79 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  spriteVisibleRegs_80 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  spriteVisibleRegs_81 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  spriteVisibleRegs_82 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  spriteVisibleRegs_83 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  spriteVisibleRegs_84 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  spriteVisibleRegs_85 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  spriteVisibleRegs_86 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  spriteVisibleRegs_87 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  spriteVisibleRegs_88 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  spriteVisibleRegs_89 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  spriteVisibleRegs_90 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  spriteVisibleRegs_91 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  spriteVisibleRegs_92 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  spriteVisibleRegs_93 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  spriteVisibleRegs_94 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  spriteVisibleRegs_95 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  spriteVisibleRegs_96 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  spriteVisibleRegs_97 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  spriteVisibleRegs_98 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  spriteVisibleRegs_99 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  spriteScaleTypeRegs_0 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  spriteScaleTypeRegs_1 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  spriteScaleTypeRegs_2 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  spriteScaleTypeRegs_3 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  spriteScaleTypeRegs_4 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  spriteScaleTypeRegs_5 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  spriteScaleTypeRegs_6 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  spriteScaleTypeRegs_7 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  spriteScaleTypeRegs_8 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  spriteScaleTypeRegs_9 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  initializePositions = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  sprite58ScaleUpHorizontal = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  sprite58ScaleUpVertical = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  sprite59ScaleUpHorizontal = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  sprite59ScaleUpVertical = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  sprite60ScaleUpHorizontal = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  sprite60ScaleUpVertical = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  viewBoxXReg = _RAND_229[9:0];
  _RAND_230 = {1{`RANDOM}};
  viewBoxYReg = _RAND_230[8:0];
  _RAND_231 = {1{`RANDOM}};
  lvlReg = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  livesReg = _RAND_232[2:0];
  _RAND_233 = {1{`RANDOM}};
  extraLifeCnt = _RAND_233[9:0];
  _RAND_234 = {1{`RANDOM}};
  gameOverReturnPressed = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  spawnDelayCounter = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  nextSpriteToSpawn = _RAND_236[5:0];
  _RAND_237 = {1{`RANDOM}};
  starCnt = _RAND_237[9:0];
  _RAND_238 = {1{`RANDOM}};
  collisionDetected = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  blinkCounter = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  blinkTimes = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  isBlinking = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  spriteXRegs_58_REG = _RAND_242[10:0];
  _RAND_243 = {1{`RANDOM}};
  spriteYRegs_58_REG = _RAND_243[9:0];
  _RAND_244 = {1{`RANDOM}};
  spriteXRegs_59_REG = _RAND_244[10:0];
  _RAND_245 = {1{`RANDOM}};
  spriteYRegs_59_REG = _RAND_245[9:0];
  _RAND_246 = {1{`RANDOM}};
  spriteXRegs_60_REG = _RAND_246[10:0];
  _RAND_247 = {1{`RANDOM}};
  spriteYRegs_60_REG = _RAND_247[9:0];
  _RAND_248 = {1{`RANDOM}};
  spriteXRegs_58_REG_1 = _RAND_248[10:0];
  _RAND_249 = {1{`RANDOM}};
  spriteYRegs_58_REG_1 = _RAND_249[9:0];
  _RAND_250 = {1{`RANDOM}};
  spriteXRegs_59_REG_1 = _RAND_250[10:0];
  _RAND_251 = {1{`RANDOM}};
  spriteYRegs_59_REG_1 = _RAND_251[9:0];
  _RAND_252 = {1{`RANDOM}};
  spriteXRegs_60_REG_1 = _RAND_252[10:0];
  _RAND_253 = {1{`RANDOM}};
  spriteYRegs_60_REG_1 = _RAND_253[9:0];
  _RAND_254 = {1{`RANDOM}};
  spriteXRegs_58_REG_2 = _RAND_254[10:0];
  _RAND_255 = {1{`RANDOM}};
  spriteYRegs_58_REG_2 = _RAND_255[9:0];
  _RAND_256 = {1{`RANDOM}};
  spriteXRegs_59_REG_2 = _RAND_256[10:0];
  _RAND_257 = {1{`RANDOM}};
  spriteYRegs_59_REG_2 = _RAND_257[9:0];
  _RAND_258 = {1{`RANDOM}};
  spriteXRegs_60_REG_2 = _RAND_258[10:0];
  _RAND_259 = {1{`RANDOM}};
  spriteYRegs_60_REG_2 = _RAND_259[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GameTop(
  input        clock,
  input        reset,
  input        io_btnC, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnU, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnL, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnR, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnD, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaRed, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaBlue, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaGreen, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_Hsync, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_Vsync, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_missingFrameError, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_viewBoxOutOfRangeError // @[\\src\\main\\scala\\GameTop.scala 14:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  graphicEngineVGA_clock; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_reset; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_46; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_47; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_48; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_49; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_50; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_51; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_52; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_53; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_54; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_55; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_56; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_57; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_61; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_62; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_63; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_46; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_47; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_48; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_49; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_50; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_51; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_52; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_53; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_54; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_55; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_56; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_57; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_61; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_62; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_63; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_46; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_47; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_48; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_49; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_50; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_51; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_52; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_53; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_54; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_55; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_56; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_57; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_61; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_62; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_63; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_64; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_65; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_66; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_67; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_68; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_69; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_70; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_71; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_72; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_73; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_74; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_75; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_76; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_77; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_78; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_79; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_80; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_81; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_82; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_83; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_84; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_85; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_86; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_87; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_88; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_89; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_90; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_91; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_92; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_93; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_94; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_95; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_96; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_97; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_98; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_99; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [8:0] graphicEngineVGA_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_missingFrameError; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaRed; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaBlue; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaGreen; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Hsync; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Vsync; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  soundEngine_clock; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  soundEngine_reset; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  gameLogic_clock; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_reset; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnC; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnU; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnL; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnR; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnD; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_46; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_47; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_48; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_49; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_50; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_51; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_52; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_53; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_54; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_55; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_56; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_57; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_61; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_62; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_63; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_46; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_47; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_48; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_49; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_50; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_51; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_52; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_53; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_54; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_55; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_56; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_57; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_61; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_62; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_63; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_46; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_47; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_48; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_49; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_50; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_51; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_52; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_53; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_54; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_55; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_56; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_57; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_61; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_62; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_63; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_64; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_65; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_66; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_67; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_68; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_69; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_70; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_71; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_72; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_73; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_74; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_75; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_76; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_77; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_78; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_79; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_80; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_81; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_82; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_83; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_84; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_85; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_86; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_87; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_88; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_89; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_90; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_91; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_92; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_93; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_94; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_95; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_96; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_97; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_98; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_99; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [8:0] gameLogic_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  reg [20:0] debounceCounter; // @[\\src\\main\\scala\\GameTop.scala 68:32]
  wire  debounceSampleEn = debounceCounter == 21'h1e847f; // @[\\src\\main\\scala\\GameTop.scala 70:24]
  wire [20:0] _debounceCounter_T_1 = debounceCounter + 21'h1; // @[\\src\\main\\scala\\GameTop.scala 74:40]
  reg [21:0] resetReleaseCounter; // @[\\src\\main\\scala\\GameTop.scala 81:36]
  wire [21:0] _resetReleaseCounter_T_1 = resetReleaseCounter + 22'h1; // @[\\src\\main\\scala\\GameTop.scala 87:48]
  reg  btnCState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnCState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnCState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnCState; // @[\\src\\main\\scala\\GameTop.scala 93:28]
  reg  btnUState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState; // @[\\src\\main\\scala\\GameTop.scala 94:28]
  reg  btnLState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState; // @[\\src\\main\\scala\\GameTop.scala 95:28]
  reg  btnRState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState; // @[\\src\\main\\scala\\GameTop.scala 96:28]
  reg  btnDState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState; // @[\\src\\main\\scala\\GameTop.scala 97:28]
  GraphicEngineVGA graphicEngineVGA ( // @[\\src\\main\\scala\\GameTop.scala 46:32]
    .clock(graphicEngineVGA_clock),
    .reset(graphicEngineVGA_reset),
    .io_spriteXPosition_3(graphicEngineVGA_io_spriteXPosition_3),
    .io_spriteXPosition_7(graphicEngineVGA_io_spriteXPosition_7),
    .io_spriteXPosition_8(graphicEngineVGA_io_spriteXPosition_8),
    .io_spriteXPosition_9(graphicEngineVGA_io_spriteXPosition_9),
    .io_spriteXPosition_10(graphicEngineVGA_io_spriteXPosition_10),
    .io_spriteXPosition_11(graphicEngineVGA_io_spriteXPosition_11),
    .io_spriteXPosition_12(graphicEngineVGA_io_spriteXPosition_12),
    .io_spriteXPosition_13(graphicEngineVGA_io_spriteXPosition_13),
    .io_spriteXPosition_14(graphicEngineVGA_io_spriteXPosition_14),
    .io_spriteXPosition_16(graphicEngineVGA_io_spriteXPosition_16),
    .io_spriteXPosition_17(graphicEngineVGA_io_spriteXPosition_17),
    .io_spriteXPosition_18(graphicEngineVGA_io_spriteXPosition_18),
    .io_spriteXPosition_19(graphicEngineVGA_io_spriteXPosition_19),
    .io_spriteXPosition_20(graphicEngineVGA_io_spriteXPosition_20),
    .io_spriteXPosition_21(graphicEngineVGA_io_spriteXPosition_21),
    .io_spriteXPosition_22(graphicEngineVGA_io_spriteXPosition_22),
    .io_spriteXPosition_23(graphicEngineVGA_io_spriteXPosition_23),
    .io_spriteXPosition_24(graphicEngineVGA_io_spriteXPosition_24),
    .io_spriteXPosition_25(graphicEngineVGA_io_spriteXPosition_25),
    .io_spriteXPosition_26(graphicEngineVGA_io_spriteXPosition_26),
    .io_spriteXPosition_27(graphicEngineVGA_io_spriteXPosition_27),
    .io_spriteXPosition_28(graphicEngineVGA_io_spriteXPosition_28),
    .io_spriteXPosition_29(graphicEngineVGA_io_spriteXPosition_29),
    .io_spriteXPosition_30(graphicEngineVGA_io_spriteXPosition_30),
    .io_spriteXPosition_31(graphicEngineVGA_io_spriteXPosition_31),
    .io_spriteXPosition_32(graphicEngineVGA_io_spriteXPosition_32),
    .io_spriteXPosition_33(graphicEngineVGA_io_spriteXPosition_33),
    .io_spriteXPosition_34(graphicEngineVGA_io_spriteXPosition_34),
    .io_spriteXPosition_35(graphicEngineVGA_io_spriteXPosition_35),
    .io_spriteXPosition_36(graphicEngineVGA_io_spriteXPosition_36),
    .io_spriteXPosition_37(graphicEngineVGA_io_spriteXPosition_37),
    .io_spriteXPosition_38(graphicEngineVGA_io_spriteXPosition_38),
    .io_spriteXPosition_39(graphicEngineVGA_io_spriteXPosition_39),
    .io_spriteXPosition_40(graphicEngineVGA_io_spriteXPosition_40),
    .io_spriteXPosition_41(graphicEngineVGA_io_spriteXPosition_41),
    .io_spriteXPosition_42(graphicEngineVGA_io_spriteXPosition_42),
    .io_spriteXPosition_43(graphicEngineVGA_io_spriteXPosition_43),
    .io_spriteXPosition_44(graphicEngineVGA_io_spriteXPosition_44),
    .io_spriteXPosition_45(graphicEngineVGA_io_spriteXPosition_45),
    .io_spriteXPosition_46(graphicEngineVGA_io_spriteXPosition_46),
    .io_spriteXPosition_47(graphicEngineVGA_io_spriteXPosition_47),
    .io_spriteXPosition_48(graphicEngineVGA_io_spriteXPosition_48),
    .io_spriteXPosition_49(graphicEngineVGA_io_spriteXPosition_49),
    .io_spriteXPosition_50(graphicEngineVGA_io_spriteXPosition_50),
    .io_spriteXPosition_51(graphicEngineVGA_io_spriteXPosition_51),
    .io_spriteXPosition_52(graphicEngineVGA_io_spriteXPosition_52),
    .io_spriteXPosition_53(graphicEngineVGA_io_spriteXPosition_53),
    .io_spriteXPosition_54(graphicEngineVGA_io_spriteXPosition_54),
    .io_spriteXPosition_55(graphicEngineVGA_io_spriteXPosition_55),
    .io_spriteXPosition_56(graphicEngineVGA_io_spriteXPosition_56),
    .io_spriteXPosition_57(graphicEngineVGA_io_spriteXPosition_57),
    .io_spriteXPosition_58(graphicEngineVGA_io_spriteXPosition_58),
    .io_spriteXPosition_59(graphicEngineVGA_io_spriteXPosition_59),
    .io_spriteXPosition_60(graphicEngineVGA_io_spriteXPosition_60),
    .io_spriteXPosition_61(graphicEngineVGA_io_spriteXPosition_61),
    .io_spriteXPosition_62(graphicEngineVGA_io_spriteXPosition_62),
    .io_spriteXPosition_63(graphicEngineVGA_io_spriteXPosition_63),
    .io_spriteYPosition_3(graphicEngineVGA_io_spriteYPosition_3),
    .io_spriteYPosition_7(graphicEngineVGA_io_spriteYPosition_7),
    .io_spriteYPosition_8(graphicEngineVGA_io_spriteYPosition_8),
    .io_spriteYPosition_9(graphicEngineVGA_io_spriteYPosition_9),
    .io_spriteYPosition_10(graphicEngineVGA_io_spriteYPosition_10),
    .io_spriteYPosition_11(graphicEngineVGA_io_spriteYPosition_11),
    .io_spriteYPosition_12(graphicEngineVGA_io_spriteYPosition_12),
    .io_spriteYPosition_13(graphicEngineVGA_io_spriteYPosition_13),
    .io_spriteYPosition_14(graphicEngineVGA_io_spriteYPosition_14),
    .io_spriteYPosition_16(graphicEngineVGA_io_spriteYPosition_16),
    .io_spriteYPosition_17(graphicEngineVGA_io_spriteYPosition_17),
    .io_spriteYPosition_18(graphicEngineVGA_io_spriteYPosition_18),
    .io_spriteYPosition_19(graphicEngineVGA_io_spriteYPosition_19),
    .io_spriteYPosition_20(graphicEngineVGA_io_spriteYPosition_20),
    .io_spriteYPosition_21(graphicEngineVGA_io_spriteYPosition_21),
    .io_spriteYPosition_22(graphicEngineVGA_io_spriteYPosition_22),
    .io_spriteYPosition_23(graphicEngineVGA_io_spriteYPosition_23),
    .io_spriteYPosition_24(graphicEngineVGA_io_spriteYPosition_24),
    .io_spriteYPosition_25(graphicEngineVGA_io_spriteYPosition_25),
    .io_spriteYPosition_26(graphicEngineVGA_io_spriteYPosition_26),
    .io_spriteYPosition_27(graphicEngineVGA_io_spriteYPosition_27),
    .io_spriteYPosition_28(graphicEngineVGA_io_spriteYPosition_28),
    .io_spriteYPosition_29(graphicEngineVGA_io_spriteYPosition_29),
    .io_spriteYPosition_30(graphicEngineVGA_io_spriteYPosition_30),
    .io_spriteYPosition_31(graphicEngineVGA_io_spriteYPosition_31),
    .io_spriteYPosition_32(graphicEngineVGA_io_spriteYPosition_32),
    .io_spriteYPosition_33(graphicEngineVGA_io_spriteYPosition_33),
    .io_spriteYPosition_34(graphicEngineVGA_io_spriteYPosition_34),
    .io_spriteYPosition_35(graphicEngineVGA_io_spriteYPosition_35),
    .io_spriteYPosition_36(graphicEngineVGA_io_spriteYPosition_36),
    .io_spriteYPosition_37(graphicEngineVGA_io_spriteYPosition_37),
    .io_spriteYPosition_38(graphicEngineVGA_io_spriteYPosition_38),
    .io_spriteYPosition_39(graphicEngineVGA_io_spriteYPosition_39),
    .io_spriteYPosition_40(graphicEngineVGA_io_spriteYPosition_40),
    .io_spriteYPosition_41(graphicEngineVGA_io_spriteYPosition_41),
    .io_spriteYPosition_42(graphicEngineVGA_io_spriteYPosition_42),
    .io_spriteYPosition_43(graphicEngineVGA_io_spriteYPosition_43),
    .io_spriteYPosition_44(graphicEngineVGA_io_spriteYPosition_44),
    .io_spriteYPosition_45(graphicEngineVGA_io_spriteYPosition_45),
    .io_spriteYPosition_46(graphicEngineVGA_io_spriteYPosition_46),
    .io_spriteYPosition_47(graphicEngineVGA_io_spriteYPosition_47),
    .io_spriteYPosition_48(graphicEngineVGA_io_spriteYPosition_48),
    .io_spriteYPosition_49(graphicEngineVGA_io_spriteYPosition_49),
    .io_spriteYPosition_50(graphicEngineVGA_io_spriteYPosition_50),
    .io_spriteYPosition_51(graphicEngineVGA_io_spriteYPosition_51),
    .io_spriteYPosition_52(graphicEngineVGA_io_spriteYPosition_52),
    .io_spriteYPosition_53(graphicEngineVGA_io_spriteYPosition_53),
    .io_spriteYPosition_54(graphicEngineVGA_io_spriteYPosition_54),
    .io_spriteYPosition_55(graphicEngineVGA_io_spriteYPosition_55),
    .io_spriteYPosition_56(graphicEngineVGA_io_spriteYPosition_56),
    .io_spriteYPosition_57(graphicEngineVGA_io_spriteYPosition_57),
    .io_spriteYPosition_58(graphicEngineVGA_io_spriteYPosition_58),
    .io_spriteYPosition_59(graphicEngineVGA_io_spriteYPosition_59),
    .io_spriteYPosition_60(graphicEngineVGA_io_spriteYPosition_60),
    .io_spriteYPosition_61(graphicEngineVGA_io_spriteYPosition_61),
    .io_spriteYPosition_62(graphicEngineVGA_io_spriteYPosition_62),
    .io_spriteYPosition_63(graphicEngineVGA_io_spriteYPosition_63),
    .io_spriteVisible_3(graphicEngineVGA_io_spriteVisible_3),
    .io_spriteVisible_4(graphicEngineVGA_io_spriteVisible_4),
    .io_spriteVisible_5(graphicEngineVGA_io_spriteVisible_5),
    .io_spriteVisible_6(graphicEngineVGA_io_spriteVisible_6),
    .io_spriteVisible_7(graphicEngineVGA_io_spriteVisible_7),
    .io_spriteVisible_8(graphicEngineVGA_io_spriteVisible_8),
    .io_spriteVisible_9(graphicEngineVGA_io_spriteVisible_9),
    .io_spriteVisible_10(graphicEngineVGA_io_spriteVisible_10),
    .io_spriteVisible_11(graphicEngineVGA_io_spriteVisible_11),
    .io_spriteVisible_12(graphicEngineVGA_io_spriteVisible_12),
    .io_spriteVisible_13(graphicEngineVGA_io_spriteVisible_13),
    .io_spriteVisible_14(graphicEngineVGA_io_spriteVisible_14),
    .io_spriteVisible_15(graphicEngineVGA_io_spriteVisible_15),
    .io_spriteVisible_16(graphicEngineVGA_io_spriteVisible_16),
    .io_spriteVisible_17(graphicEngineVGA_io_spriteVisible_17),
    .io_spriteVisible_18(graphicEngineVGA_io_spriteVisible_18),
    .io_spriteVisible_19(graphicEngineVGA_io_spriteVisible_19),
    .io_spriteVisible_20(graphicEngineVGA_io_spriteVisible_20),
    .io_spriteVisible_21(graphicEngineVGA_io_spriteVisible_21),
    .io_spriteVisible_22(graphicEngineVGA_io_spriteVisible_22),
    .io_spriteVisible_23(graphicEngineVGA_io_spriteVisible_23),
    .io_spriteVisible_24(graphicEngineVGA_io_spriteVisible_24),
    .io_spriteVisible_25(graphicEngineVGA_io_spriteVisible_25),
    .io_spriteVisible_26(graphicEngineVGA_io_spriteVisible_26),
    .io_spriteVisible_27(graphicEngineVGA_io_spriteVisible_27),
    .io_spriteVisible_28(graphicEngineVGA_io_spriteVisible_28),
    .io_spriteVisible_29(graphicEngineVGA_io_spriteVisible_29),
    .io_spriteVisible_30(graphicEngineVGA_io_spriteVisible_30),
    .io_spriteVisible_31(graphicEngineVGA_io_spriteVisible_31),
    .io_spriteVisible_32(graphicEngineVGA_io_spriteVisible_32),
    .io_spriteVisible_33(graphicEngineVGA_io_spriteVisible_33),
    .io_spriteVisible_34(graphicEngineVGA_io_spriteVisible_34),
    .io_spriteVisible_35(graphicEngineVGA_io_spriteVisible_35),
    .io_spriteVisible_36(graphicEngineVGA_io_spriteVisible_36),
    .io_spriteVisible_37(graphicEngineVGA_io_spriteVisible_37),
    .io_spriteVisible_38(graphicEngineVGA_io_spriteVisible_38),
    .io_spriteVisible_39(graphicEngineVGA_io_spriteVisible_39),
    .io_spriteVisible_40(graphicEngineVGA_io_spriteVisible_40),
    .io_spriteVisible_41(graphicEngineVGA_io_spriteVisible_41),
    .io_spriteVisible_42(graphicEngineVGA_io_spriteVisible_42),
    .io_spriteVisible_43(graphicEngineVGA_io_spriteVisible_43),
    .io_spriteVisible_44(graphicEngineVGA_io_spriteVisible_44),
    .io_spriteVisible_45(graphicEngineVGA_io_spriteVisible_45),
    .io_spriteVisible_46(graphicEngineVGA_io_spriteVisible_46),
    .io_spriteVisible_47(graphicEngineVGA_io_spriteVisible_47),
    .io_spriteVisible_48(graphicEngineVGA_io_spriteVisible_48),
    .io_spriteVisible_49(graphicEngineVGA_io_spriteVisible_49),
    .io_spriteVisible_50(graphicEngineVGA_io_spriteVisible_50),
    .io_spriteVisible_51(graphicEngineVGA_io_spriteVisible_51),
    .io_spriteVisible_52(graphicEngineVGA_io_spriteVisible_52),
    .io_spriteVisible_53(graphicEngineVGA_io_spriteVisible_53),
    .io_spriteVisible_54(graphicEngineVGA_io_spriteVisible_54),
    .io_spriteVisible_55(graphicEngineVGA_io_spriteVisible_55),
    .io_spriteVisible_56(graphicEngineVGA_io_spriteVisible_56),
    .io_spriteVisible_57(graphicEngineVGA_io_spriteVisible_57),
    .io_spriteVisible_58(graphicEngineVGA_io_spriteVisible_58),
    .io_spriteVisible_59(graphicEngineVGA_io_spriteVisible_59),
    .io_spriteVisible_60(graphicEngineVGA_io_spriteVisible_60),
    .io_spriteVisible_61(graphicEngineVGA_io_spriteVisible_61),
    .io_spriteVisible_62(graphicEngineVGA_io_spriteVisible_62),
    .io_spriteVisible_63(graphicEngineVGA_io_spriteVisible_63),
    .io_spriteVisible_64(graphicEngineVGA_io_spriteVisible_64),
    .io_spriteVisible_65(graphicEngineVGA_io_spriteVisible_65),
    .io_spriteVisible_66(graphicEngineVGA_io_spriteVisible_66),
    .io_spriteVisible_67(graphicEngineVGA_io_spriteVisible_67),
    .io_spriteVisible_68(graphicEngineVGA_io_spriteVisible_68),
    .io_spriteVisible_69(graphicEngineVGA_io_spriteVisible_69),
    .io_spriteVisible_70(graphicEngineVGA_io_spriteVisible_70),
    .io_spriteVisible_71(graphicEngineVGA_io_spriteVisible_71),
    .io_spriteVisible_72(graphicEngineVGA_io_spriteVisible_72),
    .io_spriteVisible_73(graphicEngineVGA_io_spriteVisible_73),
    .io_spriteVisible_74(graphicEngineVGA_io_spriteVisible_74),
    .io_spriteVisible_75(graphicEngineVGA_io_spriteVisible_75),
    .io_spriteVisible_76(graphicEngineVGA_io_spriteVisible_76),
    .io_spriteVisible_77(graphicEngineVGA_io_spriteVisible_77),
    .io_spriteVisible_78(graphicEngineVGA_io_spriteVisible_78),
    .io_spriteVisible_79(graphicEngineVGA_io_spriteVisible_79),
    .io_spriteVisible_80(graphicEngineVGA_io_spriteVisible_80),
    .io_spriteVisible_81(graphicEngineVGA_io_spriteVisible_81),
    .io_spriteVisible_82(graphicEngineVGA_io_spriteVisible_82),
    .io_spriteVisible_83(graphicEngineVGA_io_spriteVisible_83),
    .io_spriteVisible_84(graphicEngineVGA_io_spriteVisible_84),
    .io_spriteVisible_85(graphicEngineVGA_io_spriteVisible_85),
    .io_spriteVisible_86(graphicEngineVGA_io_spriteVisible_86),
    .io_spriteVisible_87(graphicEngineVGA_io_spriteVisible_87),
    .io_spriteVisible_88(graphicEngineVGA_io_spriteVisible_88),
    .io_spriteVisible_89(graphicEngineVGA_io_spriteVisible_89),
    .io_spriteVisible_90(graphicEngineVGA_io_spriteVisible_90),
    .io_spriteVisible_91(graphicEngineVGA_io_spriteVisible_91),
    .io_spriteVisible_92(graphicEngineVGA_io_spriteVisible_92),
    .io_spriteVisible_93(graphicEngineVGA_io_spriteVisible_93),
    .io_spriteVisible_94(graphicEngineVGA_io_spriteVisible_94),
    .io_spriteVisible_95(graphicEngineVGA_io_spriteVisible_95),
    .io_spriteVisible_96(graphicEngineVGA_io_spriteVisible_96),
    .io_spriteVisible_97(graphicEngineVGA_io_spriteVisible_97),
    .io_spriteVisible_98(graphicEngineVGA_io_spriteVisible_98),
    .io_spriteVisible_99(graphicEngineVGA_io_spriteVisible_99),
    .io_spriteScaleUpHorizontal_16(graphicEngineVGA_io_spriteScaleUpHorizontal_16),
    .io_spriteScaleUpHorizontal_17(graphicEngineVGA_io_spriteScaleUpHorizontal_17),
    .io_spriteScaleUpHorizontal_18(graphicEngineVGA_io_spriteScaleUpHorizontal_18),
    .io_spriteScaleUpHorizontal_19(graphicEngineVGA_io_spriteScaleUpHorizontal_19),
    .io_spriteScaleUpHorizontal_20(graphicEngineVGA_io_spriteScaleUpHorizontal_20),
    .io_spriteScaleUpHorizontal_21(graphicEngineVGA_io_spriteScaleUpHorizontal_21),
    .io_spriteScaleUpHorizontal_22(graphicEngineVGA_io_spriteScaleUpHorizontal_22),
    .io_spriteScaleUpHorizontal_23(graphicEngineVGA_io_spriteScaleUpHorizontal_23),
    .io_spriteScaleUpHorizontal_24(graphicEngineVGA_io_spriteScaleUpHorizontal_24),
    .io_spriteScaleUpHorizontal_25(graphicEngineVGA_io_spriteScaleUpHorizontal_25),
    .io_spriteScaleUpHorizontal_26(graphicEngineVGA_io_spriteScaleUpHorizontal_26),
    .io_spriteScaleUpHorizontal_27(graphicEngineVGA_io_spriteScaleUpHorizontal_27),
    .io_spriteScaleUpHorizontal_28(graphicEngineVGA_io_spriteScaleUpHorizontal_28),
    .io_spriteScaleUpHorizontal_29(graphicEngineVGA_io_spriteScaleUpHorizontal_29),
    .io_spriteScaleUpHorizontal_30(graphicEngineVGA_io_spriteScaleUpHorizontal_30),
    .io_spriteScaleUpHorizontal_31(graphicEngineVGA_io_spriteScaleUpHorizontal_31),
    .io_spriteScaleUpHorizontal_32(graphicEngineVGA_io_spriteScaleUpHorizontal_32),
    .io_spriteScaleUpHorizontal_33(graphicEngineVGA_io_spriteScaleUpHorizontal_33),
    .io_spriteScaleUpHorizontal_34(graphicEngineVGA_io_spriteScaleUpHorizontal_34),
    .io_spriteScaleUpHorizontal_35(graphicEngineVGA_io_spriteScaleUpHorizontal_35),
    .io_spriteScaleUpHorizontal_36(graphicEngineVGA_io_spriteScaleUpHorizontal_36),
    .io_spriteScaleUpHorizontal_37(graphicEngineVGA_io_spriteScaleUpHorizontal_37),
    .io_spriteScaleUpHorizontal_38(graphicEngineVGA_io_spriteScaleUpHorizontal_38),
    .io_spriteScaleUpHorizontal_39(graphicEngineVGA_io_spriteScaleUpHorizontal_39),
    .io_spriteScaleUpHorizontal_40(graphicEngineVGA_io_spriteScaleUpHorizontal_40),
    .io_spriteScaleUpHorizontal_41(graphicEngineVGA_io_spriteScaleUpHorizontal_41),
    .io_spriteScaleUpHorizontal_42(graphicEngineVGA_io_spriteScaleUpHorizontal_42),
    .io_spriteScaleUpHorizontal_43(graphicEngineVGA_io_spriteScaleUpHorizontal_43),
    .io_spriteScaleUpHorizontal_44(graphicEngineVGA_io_spriteScaleUpHorizontal_44),
    .io_spriteScaleUpHorizontal_45(graphicEngineVGA_io_spriteScaleUpHorizontal_45),
    .io_spriteScaleUpHorizontal_58(graphicEngineVGA_io_spriteScaleUpHorizontal_58),
    .io_spriteScaleUpHorizontal_59(graphicEngineVGA_io_spriteScaleUpHorizontal_59),
    .io_spriteScaleUpHorizontal_60(graphicEngineVGA_io_spriteScaleUpHorizontal_60),
    .io_spriteScaleUpVertical_16(graphicEngineVGA_io_spriteScaleUpVertical_16),
    .io_spriteScaleUpVertical_17(graphicEngineVGA_io_spriteScaleUpVertical_17),
    .io_spriteScaleUpVertical_18(graphicEngineVGA_io_spriteScaleUpVertical_18),
    .io_spriteScaleUpVertical_19(graphicEngineVGA_io_spriteScaleUpVertical_19),
    .io_spriteScaleUpVertical_20(graphicEngineVGA_io_spriteScaleUpVertical_20),
    .io_spriteScaleUpVertical_21(graphicEngineVGA_io_spriteScaleUpVertical_21),
    .io_spriteScaleUpVertical_22(graphicEngineVGA_io_spriteScaleUpVertical_22),
    .io_spriteScaleUpVertical_23(graphicEngineVGA_io_spriteScaleUpVertical_23),
    .io_spriteScaleUpVertical_24(graphicEngineVGA_io_spriteScaleUpVertical_24),
    .io_spriteScaleUpVertical_25(graphicEngineVGA_io_spriteScaleUpVertical_25),
    .io_spriteScaleUpVertical_26(graphicEngineVGA_io_spriteScaleUpVertical_26),
    .io_spriteScaleUpVertical_27(graphicEngineVGA_io_spriteScaleUpVertical_27),
    .io_spriteScaleUpVertical_28(graphicEngineVGA_io_spriteScaleUpVertical_28),
    .io_spriteScaleUpVertical_29(graphicEngineVGA_io_spriteScaleUpVertical_29),
    .io_spriteScaleUpVertical_30(graphicEngineVGA_io_spriteScaleUpVertical_30),
    .io_spriteScaleUpVertical_31(graphicEngineVGA_io_spriteScaleUpVertical_31),
    .io_spriteScaleUpVertical_32(graphicEngineVGA_io_spriteScaleUpVertical_32),
    .io_spriteScaleUpVertical_33(graphicEngineVGA_io_spriteScaleUpVertical_33),
    .io_spriteScaleUpVertical_34(graphicEngineVGA_io_spriteScaleUpVertical_34),
    .io_spriteScaleUpVertical_35(graphicEngineVGA_io_spriteScaleUpVertical_35),
    .io_spriteScaleUpVertical_36(graphicEngineVGA_io_spriteScaleUpVertical_36),
    .io_spriteScaleUpVertical_37(graphicEngineVGA_io_spriteScaleUpVertical_37),
    .io_spriteScaleUpVertical_38(graphicEngineVGA_io_spriteScaleUpVertical_38),
    .io_spriteScaleUpVertical_39(graphicEngineVGA_io_spriteScaleUpVertical_39),
    .io_spriteScaleUpVertical_40(graphicEngineVGA_io_spriteScaleUpVertical_40),
    .io_spriteScaleUpVertical_41(graphicEngineVGA_io_spriteScaleUpVertical_41),
    .io_spriteScaleUpVertical_42(graphicEngineVGA_io_spriteScaleUpVertical_42),
    .io_spriteScaleUpVertical_43(graphicEngineVGA_io_spriteScaleUpVertical_43),
    .io_spriteScaleUpVertical_44(graphicEngineVGA_io_spriteScaleUpVertical_44),
    .io_spriteScaleUpVertical_45(graphicEngineVGA_io_spriteScaleUpVertical_45),
    .io_spriteScaleUpVertical_58(graphicEngineVGA_io_spriteScaleUpVertical_58),
    .io_spriteScaleUpVertical_59(graphicEngineVGA_io_spriteScaleUpVertical_59),
    .io_spriteScaleUpVertical_60(graphicEngineVGA_io_spriteScaleUpVertical_60),
    .io_viewBoxX(graphicEngineVGA_io_viewBoxX),
    .io_viewBoxY(graphicEngineVGA_io_viewBoxY),
    .io_newFrame(graphicEngineVGA_io_newFrame),
    .io_frameUpdateDone(graphicEngineVGA_io_frameUpdateDone),
    .io_missingFrameError(graphicEngineVGA_io_missingFrameError),
    .io_viewBoxOutOfRangeError(graphicEngineVGA_io_viewBoxOutOfRangeError),
    .io_vgaRed(graphicEngineVGA_io_vgaRed),
    .io_vgaBlue(graphicEngineVGA_io_vgaBlue),
    .io_vgaGreen(graphicEngineVGA_io_vgaGreen),
    .io_Hsync(graphicEngineVGA_io_Hsync),
    .io_Vsync(graphicEngineVGA_io_Vsync)
  );
  SoundEngine soundEngine ( // @[\\src\\main\\scala\\GameTop.scala 49:27]
    .clock(soundEngine_clock),
    .reset(soundEngine_reset)
  );
  GameLogic gameLogic ( // @[\\src\\main\\scala\\GameTop.scala 53:25]
    .clock(gameLogic_clock),
    .reset(gameLogic_reset),
    .io_btnC(gameLogic_io_btnC),
    .io_btnU(gameLogic_io_btnU),
    .io_btnL(gameLogic_io_btnL),
    .io_btnR(gameLogic_io_btnR),
    .io_btnD(gameLogic_io_btnD),
    .io_spriteXPosition_3(gameLogic_io_spriteXPosition_3),
    .io_spriteXPosition_7(gameLogic_io_spriteXPosition_7),
    .io_spriteXPosition_8(gameLogic_io_spriteXPosition_8),
    .io_spriteXPosition_9(gameLogic_io_spriteXPosition_9),
    .io_spriteXPosition_10(gameLogic_io_spriteXPosition_10),
    .io_spriteXPosition_11(gameLogic_io_spriteXPosition_11),
    .io_spriteXPosition_12(gameLogic_io_spriteXPosition_12),
    .io_spriteXPosition_13(gameLogic_io_spriteXPosition_13),
    .io_spriteXPosition_14(gameLogic_io_spriteXPosition_14),
    .io_spriteXPosition_16(gameLogic_io_spriteXPosition_16),
    .io_spriteXPosition_17(gameLogic_io_spriteXPosition_17),
    .io_spriteXPosition_18(gameLogic_io_spriteXPosition_18),
    .io_spriteXPosition_19(gameLogic_io_spriteXPosition_19),
    .io_spriteXPosition_20(gameLogic_io_spriteXPosition_20),
    .io_spriteXPosition_21(gameLogic_io_spriteXPosition_21),
    .io_spriteXPosition_22(gameLogic_io_spriteXPosition_22),
    .io_spriteXPosition_23(gameLogic_io_spriteXPosition_23),
    .io_spriteXPosition_24(gameLogic_io_spriteXPosition_24),
    .io_spriteXPosition_25(gameLogic_io_spriteXPosition_25),
    .io_spriteXPosition_26(gameLogic_io_spriteXPosition_26),
    .io_spriteXPosition_27(gameLogic_io_spriteXPosition_27),
    .io_spriteXPosition_28(gameLogic_io_spriteXPosition_28),
    .io_spriteXPosition_29(gameLogic_io_spriteXPosition_29),
    .io_spriteXPosition_30(gameLogic_io_spriteXPosition_30),
    .io_spriteXPosition_31(gameLogic_io_spriteXPosition_31),
    .io_spriteXPosition_32(gameLogic_io_spriteXPosition_32),
    .io_spriteXPosition_33(gameLogic_io_spriteXPosition_33),
    .io_spriteXPosition_34(gameLogic_io_spriteXPosition_34),
    .io_spriteXPosition_35(gameLogic_io_spriteXPosition_35),
    .io_spriteXPosition_36(gameLogic_io_spriteXPosition_36),
    .io_spriteXPosition_37(gameLogic_io_spriteXPosition_37),
    .io_spriteXPosition_38(gameLogic_io_spriteXPosition_38),
    .io_spriteXPosition_39(gameLogic_io_spriteXPosition_39),
    .io_spriteXPosition_40(gameLogic_io_spriteXPosition_40),
    .io_spriteXPosition_41(gameLogic_io_spriteXPosition_41),
    .io_spriteXPosition_42(gameLogic_io_spriteXPosition_42),
    .io_spriteXPosition_43(gameLogic_io_spriteXPosition_43),
    .io_spriteXPosition_44(gameLogic_io_spriteXPosition_44),
    .io_spriteXPosition_45(gameLogic_io_spriteXPosition_45),
    .io_spriteXPosition_46(gameLogic_io_spriteXPosition_46),
    .io_spriteXPosition_47(gameLogic_io_spriteXPosition_47),
    .io_spriteXPosition_48(gameLogic_io_spriteXPosition_48),
    .io_spriteXPosition_49(gameLogic_io_spriteXPosition_49),
    .io_spriteXPosition_50(gameLogic_io_spriteXPosition_50),
    .io_spriteXPosition_51(gameLogic_io_spriteXPosition_51),
    .io_spriteXPosition_52(gameLogic_io_spriteXPosition_52),
    .io_spriteXPosition_53(gameLogic_io_spriteXPosition_53),
    .io_spriteXPosition_54(gameLogic_io_spriteXPosition_54),
    .io_spriteXPosition_55(gameLogic_io_spriteXPosition_55),
    .io_spriteXPosition_56(gameLogic_io_spriteXPosition_56),
    .io_spriteXPosition_57(gameLogic_io_spriteXPosition_57),
    .io_spriteXPosition_58(gameLogic_io_spriteXPosition_58),
    .io_spriteXPosition_59(gameLogic_io_spriteXPosition_59),
    .io_spriteXPosition_60(gameLogic_io_spriteXPosition_60),
    .io_spriteXPosition_61(gameLogic_io_spriteXPosition_61),
    .io_spriteXPosition_62(gameLogic_io_spriteXPosition_62),
    .io_spriteXPosition_63(gameLogic_io_spriteXPosition_63),
    .io_spriteYPosition_3(gameLogic_io_spriteYPosition_3),
    .io_spriteYPosition_7(gameLogic_io_spriteYPosition_7),
    .io_spriteYPosition_8(gameLogic_io_spriteYPosition_8),
    .io_spriteYPosition_9(gameLogic_io_spriteYPosition_9),
    .io_spriteYPosition_10(gameLogic_io_spriteYPosition_10),
    .io_spriteYPosition_11(gameLogic_io_spriteYPosition_11),
    .io_spriteYPosition_12(gameLogic_io_spriteYPosition_12),
    .io_spriteYPosition_13(gameLogic_io_spriteYPosition_13),
    .io_spriteYPosition_14(gameLogic_io_spriteYPosition_14),
    .io_spriteYPosition_16(gameLogic_io_spriteYPosition_16),
    .io_spriteYPosition_17(gameLogic_io_spriteYPosition_17),
    .io_spriteYPosition_18(gameLogic_io_spriteYPosition_18),
    .io_spriteYPosition_19(gameLogic_io_spriteYPosition_19),
    .io_spriteYPosition_20(gameLogic_io_spriteYPosition_20),
    .io_spriteYPosition_21(gameLogic_io_spriteYPosition_21),
    .io_spriteYPosition_22(gameLogic_io_spriteYPosition_22),
    .io_spriteYPosition_23(gameLogic_io_spriteYPosition_23),
    .io_spriteYPosition_24(gameLogic_io_spriteYPosition_24),
    .io_spriteYPosition_25(gameLogic_io_spriteYPosition_25),
    .io_spriteYPosition_26(gameLogic_io_spriteYPosition_26),
    .io_spriteYPosition_27(gameLogic_io_spriteYPosition_27),
    .io_spriteYPosition_28(gameLogic_io_spriteYPosition_28),
    .io_spriteYPosition_29(gameLogic_io_spriteYPosition_29),
    .io_spriteYPosition_30(gameLogic_io_spriteYPosition_30),
    .io_spriteYPosition_31(gameLogic_io_spriteYPosition_31),
    .io_spriteYPosition_32(gameLogic_io_spriteYPosition_32),
    .io_spriteYPosition_33(gameLogic_io_spriteYPosition_33),
    .io_spriteYPosition_34(gameLogic_io_spriteYPosition_34),
    .io_spriteYPosition_35(gameLogic_io_spriteYPosition_35),
    .io_spriteYPosition_36(gameLogic_io_spriteYPosition_36),
    .io_spriteYPosition_37(gameLogic_io_spriteYPosition_37),
    .io_spriteYPosition_38(gameLogic_io_spriteYPosition_38),
    .io_spriteYPosition_39(gameLogic_io_spriteYPosition_39),
    .io_spriteYPosition_40(gameLogic_io_spriteYPosition_40),
    .io_spriteYPosition_41(gameLogic_io_spriteYPosition_41),
    .io_spriteYPosition_42(gameLogic_io_spriteYPosition_42),
    .io_spriteYPosition_43(gameLogic_io_spriteYPosition_43),
    .io_spriteYPosition_44(gameLogic_io_spriteYPosition_44),
    .io_spriteYPosition_45(gameLogic_io_spriteYPosition_45),
    .io_spriteYPosition_46(gameLogic_io_spriteYPosition_46),
    .io_spriteYPosition_47(gameLogic_io_spriteYPosition_47),
    .io_spriteYPosition_48(gameLogic_io_spriteYPosition_48),
    .io_spriteYPosition_49(gameLogic_io_spriteYPosition_49),
    .io_spriteYPosition_50(gameLogic_io_spriteYPosition_50),
    .io_spriteYPosition_51(gameLogic_io_spriteYPosition_51),
    .io_spriteYPosition_52(gameLogic_io_spriteYPosition_52),
    .io_spriteYPosition_53(gameLogic_io_spriteYPosition_53),
    .io_spriteYPosition_54(gameLogic_io_spriteYPosition_54),
    .io_spriteYPosition_55(gameLogic_io_spriteYPosition_55),
    .io_spriteYPosition_56(gameLogic_io_spriteYPosition_56),
    .io_spriteYPosition_57(gameLogic_io_spriteYPosition_57),
    .io_spriteYPosition_58(gameLogic_io_spriteYPosition_58),
    .io_spriteYPosition_59(gameLogic_io_spriteYPosition_59),
    .io_spriteYPosition_60(gameLogic_io_spriteYPosition_60),
    .io_spriteYPosition_61(gameLogic_io_spriteYPosition_61),
    .io_spriteYPosition_62(gameLogic_io_spriteYPosition_62),
    .io_spriteYPosition_63(gameLogic_io_spriteYPosition_63),
    .io_spriteVisible_3(gameLogic_io_spriteVisible_3),
    .io_spriteVisible_4(gameLogic_io_spriteVisible_4),
    .io_spriteVisible_5(gameLogic_io_spriteVisible_5),
    .io_spriteVisible_6(gameLogic_io_spriteVisible_6),
    .io_spriteVisible_7(gameLogic_io_spriteVisible_7),
    .io_spriteVisible_8(gameLogic_io_spriteVisible_8),
    .io_spriteVisible_9(gameLogic_io_spriteVisible_9),
    .io_spriteVisible_10(gameLogic_io_spriteVisible_10),
    .io_spriteVisible_11(gameLogic_io_spriteVisible_11),
    .io_spriteVisible_12(gameLogic_io_spriteVisible_12),
    .io_spriteVisible_13(gameLogic_io_spriteVisible_13),
    .io_spriteVisible_14(gameLogic_io_spriteVisible_14),
    .io_spriteVisible_15(gameLogic_io_spriteVisible_15),
    .io_spriteVisible_16(gameLogic_io_spriteVisible_16),
    .io_spriteVisible_17(gameLogic_io_spriteVisible_17),
    .io_spriteVisible_18(gameLogic_io_spriteVisible_18),
    .io_spriteVisible_19(gameLogic_io_spriteVisible_19),
    .io_spriteVisible_20(gameLogic_io_spriteVisible_20),
    .io_spriteVisible_21(gameLogic_io_spriteVisible_21),
    .io_spriteVisible_22(gameLogic_io_spriteVisible_22),
    .io_spriteVisible_23(gameLogic_io_spriteVisible_23),
    .io_spriteVisible_24(gameLogic_io_spriteVisible_24),
    .io_spriteVisible_25(gameLogic_io_spriteVisible_25),
    .io_spriteVisible_26(gameLogic_io_spriteVisible_26),
    .io_spriteVisible_27(gameLogic_io_spriteVisible_27),
    .io_spriteVisible_28(gameLogic_io_spriteVisible_28),
    .io_spriteVisible_29(gameLogic_io_spriteVisible_29),
    .io_spriteVisible_30(gameLogic_io_spriteVisible_30),
    .io_spriteVisible_31(gameLogic_io_spriteVisible_31),
    .io_spriteVisible_32(gameLogic_io_spriteVisible_32),
    .io_spriteVisible_33(gameLogic_io_spriteVisible_33),
    .io_spriteVisible_34(gameLogic_io_spriteVisible_34),
    .io_spriteVisible_35(gameLogic_io_spriteVisible_35),
    .io_spriteVisible_36(gameLogic_io_spriteVisible_36),
    .io_spriteVisible_37(gameLogic_io_spriteVisible_37),
    .io_spriteVisible_38(gameLogic_io_spriteVisible_38),
    .io_spriteVisible_39(gameLogic_io_spriteVisible_39),
    .io_spriteVisible_40(gameLogic_io_spriteVisible_40),
    .io_spriteVisible_41(gameLogic_io_spriteVisible_41),
    .io_spriteVisible_42(gameLogic_io_spriteVisible_42),
    .io_spriteVisible_43(gameLogic_io_spriteVisible_43),
    .io_spriteVisible_44(gameLogic_io_spriteVisible_44),
    .io_spriteVisible_45(gameLogic_io_spriteVisible_45),
    .io_spriteVisible_46(gameLogic_io_spriteVisible_46),
    .io_spriteVisible_47(gameLogic_io_spriteVisible_47),
    .io_spriteVisible_48(gameLogic_io_spriteVisible_48),
    .io_spriteVisible_49(gameLogic_io_spriteVisible_49),
    .io_spriteVisible_50(gameLogic_io_spriteVisible_50),
    .io_spriteVisible_51(gameLogic_io_spriteVisible_51),
    .io_spriteVisible_52(gameLogic_io_spriteVisible_52),
    .io_spriteVisible_53(gameLogic_io_spriteVisible_53),
    .io_spriteVisible_54(gameLogic_io_spriteVisible_54),
    .io_spriteVisible_55(gameLogic_io_spriteVisible_55),
    .io_spriteVisible_56(gameLogic_io_spriteVisible_56),
    .io_spriteVisible_57(gameLogic_io_spriteVisible_57),
    .io_spriteVisible_58(gameLogic_io_spriteVisible_58),
    .io_spriteVisible_59(gameLogic_io_spriteVisible_59),
    .io_spriteVisible_60(gameLogic_io_spriteVisible_60),
    .io_spriteVisible_61(gameLogic_io_spriteVisible_61),
    .io_spriteVisible_62(gameLogic_io_spriteVisible_62),
    .io_spriteVisible_63(gameLogic_io_spriteVisible_63),
    .io_spriteVisible_64(gameLogic_io_spriteVisible_64),
    .io_spriteVisible_65(gameLogic_io_spriteVisible_65),
    .io_spriteVisible_66(gameLogic_io_spriteVisible_66),
    .io_spriteVisible_67(gameLogic_io_spriteVisible_67),
    .io_spriteVisible_68(gameLogic_io_spriteVisible_68),
    .io_spriteVisible_69(gameLogic_io_spriteVisible_69),
    .io_spriteVisible_70(gameLogic_io_spriteVisible_70),
    .io_spriteVisible_71(gameLogic_io_spriteVisible_71),
    .io_spriteVisible_72(gameLogic_io_spriteVisible_72),
    .io_spriteVisible_73(gameLogic_io_spriteVisible_73),
    .io_spriteVisible_74(gameLogic_io_spriteVisible_74),
    .io_spriteVisible_75(gameLogic_io_spriteVisible_75),
    .io_spriteVisible_76(gameLogic_io_spriteVisible_76),
    .io_spriteVisible_77(gameLogic_io_spriteVisible_77),
    .io_spriteVisible_78(gameLogic_io_spriteVisible_78),
    .io_spriteVisible_79(gameLogic_io_spriteVisible_79),
    .io_spriteVisible_80(gameLogic_io_spriteVisible_80),
    .io_spriteVisible_81(gameLogic_io_spriteVisible_81),
    .io_spriteVisible_82(gameLogic_io_spriteVisible_82),
    .io_spriteVisible_83(gameLogic_io_spriteVisible_83),
    .io_spriteVisible_84(gameLogic_io_spriteVisible_84),
    .io_spriteVisible_85(gameLogic_io_spriteVisible_85),
    .io_spriteVisible_86(gameLogic_io_spriteVisible_86),
    .io_spriteVisible_87(gameLogic_io_spriteVisible_87),
    .io_spriteVisible_88(gameLogic_io_spriteVisible_88),
    .io_spriteVisible_89(gameLogic_io_spriteVisible_89),
    .io_spriteVisible_90(gameLogic_io_spriteVisible_90),
    .io_spriteVisible_91(gameLogic_io_spriteVisible_91),
    .io_spriteVisible_92(gameLogic_io_spriteVisible_92),
    .io_spriteVisible_93(gameLogic_io_spriteVisible_93),
    .io_spriteVisible_94(gameLogic_io_spriteVisible_94),
    .io_spriteVisible_95(gameLogic_io_spriteVisible_95),
    .io_spriteVisible_96(gameLogic_io_spriteVisible_96),
    .io_spriteVisible_97(gameLogic_io_spriteVisible_97),
    .io_spriteVisible_98(gameLogic_io_spriteVisible_98),
    .io_spriteVisible_99(gameLogic_io_spriteVisible_99),
    .io_spriteScaleUpHorizontal_16(gameLogic_io_spriteScaleUpHorizontal_16),
    .io_spriteScaleUpHorizontal_17(gameLogic_io_spriteScaleUpHorizontal_17),
    .io_spriteScaleUpHorizontal_18(gameLogic_io_spriteScaleUpHorizontal_18),
    .io_spriteScaleUpHorizontal_19(gameLogic_io_spriteScaleUpHorizontal_19),
    .io_spriteScaleUpHorizontal_20(gameLogic_io_spriteScaleUpHorizontal_20),
    .io_spriteScaleUpHorizontal_21(gameLogic_io_spriteScaleUpHorizontal_21),
    .io_spriteScaleUpHorizontal_22(gameLogic_io_spriteScaleUpHorizontal_22),
    .io_spriteScaleUpHorizontal_23(gameLogic_io_spriteScaleUpHorizontal_23),
    .io_spriteScaleUpHorizontal_24(gameLogic_io_spriteScaleUpHorizontal_24),
    .io_spriteScaleUpHorizontal_25(gameLogic_io_spriteScaleUpHorizontal_25),
    .io_spriteScaleUpHorizontal_26(gameLogic_io_spriteScaleUpHorizontal_26),
    .io_spriteScaleUpHorizontal_27(gameLogic_io_spriteScaleUpHorizontal_27),
    .io_spriteScaleUpHorizontal_28(gameLogic_io_spriteScaleUpHorizontal_28),
    .io_spriteScaleUpHorizontal_29(gameLogic_io_spriteScaleUpHorizontal_29),
    .io_spriteScaleUpHorizontal_30(gameLogic_io_spriteScaleUpHorizontal_30),
    .io_spriteScaleUpHorizontal_31(gameLogic_io_spriteScaleUpHorizontal_31),
    .io_spriteScaleUpHorizontal_32(gameLogic_io_spriteScaleUpHorizontal_32),
    .io_spriteScaleUpHorizontal_33(gameLogic_io_spriteScaleUpHorizontal_33),
    .io_spriteScaleUpHorizontal_34(gameLogic_io_spriteScaleUpHorizontal_34),
    .io_spriteScaleUpHorizontal_35(gameLogic_io_spriteScaleUpHorizontal_35),
    .io_spriteScaleUpHorizontal_36(gameLogic_io_spriteScaleUpHorizontal_36),
    .io_spriteScaleUpHorizontal_37(gameLogic_io_spriteScaleUpHorizontal_37),
    .io_spriteScaleUpHorizontal_38(gameLogic_io_spriteScaleUpHorizontal_38),
    .io_spriteScaleUpHorizontal_39(gameLogic_io_spriteScaleUpHorizontal_39),
    .io_spriteScaleUpHorizontal_40(gameLogic_io_spriteScaleUpHorizontal_40),
    .io_spriteScaleUpHorizontal_41(gameLogic_io_spriteScaleUpHorizontal_41),
    .io_spriteScaleUpHorizontal_42(gameLogic_io_spriteScaleUpHorizontal_42),
    .io_spriteScaleUpHorizontal_43(gameLogic_io_spriteScaleUpHorizontal_43),
    .io_spriteScaleUpHorizontal_44(gameLogic_io_spriteScaleUpHorizontal_44),
    .io_spriteScaleUpHorizontal_45(gameLogic_io_spriteScaleUpHorizontal_45),
    .io_spriteScaleUpHorizontal_58(gameLogic_io_spriteScaleUpHorizontal_58),
    .io_spriteScaleUpHorizontal_59(gameLogic_io_spriteScaleUpHorizontal_59),
    .io_spriteScaleUpHorizontal_60(gameLogic_io_spriteScaleUpHorizontal_60),
    .io_spriteScaleUpVertical_16(gameLogic_io_spriteScaleUpVertical_16),
    .io_spriteScaleUpVertical_17(gameLogic_io_spriteScaleUpVertical_17),
    .io_spriteScaleUpVertical_18(gameLogic_io_spriteScaleUpVertical_18),
    .io_spriteScaleUpVertical_19(gameLogic_io_spriteScaleUpVertical_19),
    .io_spriteScaleUpVertical_20(gameLogic_io_spriteScaleUpVertical_20),
    .io_spriteScaleUpVertical_21(gameLogic_io_spriteScaleUpVertical_21),
    .io_spriteScaleUpVertical_22(gameLogic_io_spriteScaleUpVertical_22),
    .io_spriteScaleUpVertical_23(gameLogic_io_spriteScaleUpVertical_23),
    .io_spriteScaleUpVertical_24(gameLogic_io_spriteScaleUpVertical_24),
    .io_spriteScaleUpVertical_25(gameLogic_io_spriteScaleUpVertical_25),
    .io_spriteScaleUpVertical_26(gameLogic_io_spriteScaleUpVertical_26),
    .io_spriteScaleUpVertical_27(gameLogic_io_spriteScaleUpVertical_27),
    .io_spriteScaleUpVertical_28(gameLogic_io_spriteScaleUpVertical_28),
    .io_spriteScaleUpVertical_29(gameLogic_io_spriteScaleUpVertical_29),
    .io_spriteScaleUpVertical_30(gameLogic_io_spriteScaleUpVertical_30),
    .io_spriteScaleUpVertical_31(gameLogic_io_spriteScaleUpVertical_31),
    .io_spriteScaleUpVertical_32(gameLogic_io_spriteScaleUpVertical_32),
    .io_spriteScaleUpVertical_33(gameLogic_io_spriteScaleUpVertical_33),
    .io_spriteScaleUpVertical_34(gameLogic_io_spriteScaleUpVertical_34),
    .io_spriteScaleUpVertical_35(gameLogic_io_spriteScaleUpVertical_35),
    .io_spriteScaleUpVertical_36(gameLogic_io_spriteScaleUpVertical_36),
    .io_spriteScaleUpVertical_37(gameLogic_io_spriteScaleUpVertical_37),
    .io_spriteScaleUpVertical_38(gameLogic_io_spriteScaleUpVertical_38),
    .io_spriteScaleUpVertical_39(gameLogic_io_spriteScaleUpVertical_39),
    .io_spriteScaleUpVertical_40(gameLogic_io_spriteScaleUpVertical_40),
    .io_spriteScaleUpVertical_41(gameLogic_io_spriteScaleUpVertical_41),
    .io_spriteScaleUpVertical_42(gameLogic_io_spriteScaleUpVertical_42),
    .io_spriteScaleUpVertical_43(gameLogic_io_spriteScaleUpVertical_43),
    .io_spriteScaleUpVertical_44(gameLogic_io_spriteScaleUpVertical_44),
    .io_spriteScaleUpVertical_45(gameLogic_io_spriteScaleUpVertical_45),
    .io_spriteScaleUpVertical_58(gameLogic_io_spriteScaleUpVertical_58),
    .io_spriteScaleUpVertical_59(gameLogic_io_spriteScaleUpVertical_59),
    .io_spriteScaleUpVertical_60(gameLogic_io_spriteScaleUpVertical_60),
    .io_viewBoxX(gameLogic_io_viewBoxX),
    .io_viewBoxY(gameLogic_io_viewBoxY),
    .io_newFrame(gameLogic_io_newFrame),
    .io_frameUpdateDone(gameLogic_io_frameUpdateDone)
  );
  assign io_vgaRed = graphicEngineVGA_io_vgaRed; // @[\\src\\main\\scala\\GameTop.scala 105:13]
  assign io_vgaBlue = graphicEngineVGA_io_vgaBlue; // @[\\src\\main\\scala\\GameTop.scala 107:14]
  assign io_vgaGreen = graphicEngineVGA_io_vgaGreen; // @[\\src\\main\\scala\\GameTop.scala 106:15]
  assign io_Hsync = graphicEngineVGA_io_Hsync; // @[\\src\\main\\scala\\GameTop.scala 108:12]
  assign io_Vsync = graphicEngineVGA_io_Vsync; // @[\\src\\main\\scala\\GameTop.scala 109:12]
  assign io_missingFrameError = graphicEngineVGA_io_missingFrameError; // @[\\src\\main\\scala\\GameTop.scala 120:24]
  assign io_viewBoxOutOfRangeError = graphicEngineVGA_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\GameTop.scala 122:29]
  assign graphicEngineVGA_clock = clock;
  assign graphicEngineVGA_reset = resetReleaseCounter == 22'h3d08ff ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameTop.scala 83:67 84:18 86:18]
  assign graphicEngineVGA_io_spriteXPosition_3 = gameLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_7 = gameLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_8 = gameLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_9 = gameLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_10 = gameLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_11 = gameLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_12 = gameLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_13 = gameLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_14 = gameLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_16 = gameLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_17 = gameLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_18 = gameLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_19 = gameLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_20 = gameLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_21 = gameLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_22 = gameLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_23 = gameLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_24 = gameLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_25 = gameLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_26 = gameLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_27 = gameLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_28 = gameLogic_io_spriteXPosition_28; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_29 = gameLogic_io_spriteXPosition_29; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_30 = gameLogic_io_spriteXPosition_30; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_31 = gameLogic_io_spriteXPosition_31; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_32 = gameLogic_io_spriteXPosition_32; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_33 = gameLogic_io_spriteXPosition_33; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_34 = gameLogic_io_spriteXPosition_34; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_35 = gameLogic_io_spriteXPosition_35; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_36 = gameLogic_io_spriteXPosition_36; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_37 = gameLogic_io_spriteXPosition_37; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_38 = gameLogic_io_spriteXPosition_38; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_39 = gameLogic_io_spriteXPosition_39; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_40 = gameLogic_io_spriteXPosition_40; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_41 = gameLogic_io_spriteXPosition_41; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_42 = gameLogic_io_spriteXPosition_42; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_43 = gameLogic_io_spriteXPosition_43; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_44 = gameLogic_io_spriteXPosition_44; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_45 = gameLogic_io_spriteXPosition_45; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_46 = gameLogic_io_spriteXPosition_46; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_47 = gameLogic_io_spriteXPosition_47; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_48 = gameLogic_io_spriteXPosition_48; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_49 = gameLogic_io_spriteXPosition_49; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_50 = gameLogic_io_spriteXPosition_50; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_51 = gameLogic_io_spriteXPosition_51; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_52 = gameLogic_io_spriteXPosition_52; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_53 = gameLogic_io_spriteXPosition_53; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_54 = gameLogic_io_spriteXPosition_54; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_55 = gameLogic_io_spriteXPosition_55; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_56 = gameLogic_io_spriteXPosition_56; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_57 = gameLogic_io_spriteXPosition_57; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_58 = gameLogic_io_spriteXPosition_58; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_59 = gameLogic_io_spriteXPosition_59; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_60 = gameLogic_io_spriteXPosition_60; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_61 = gameLogic_io_spriteXPosition_61; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_62 = gameLogic_io_spriteXPosition_62; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_63 = gameLogic_io_spriteXPosition_63; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteYPosition_3 = gameLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_7 = gameLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_8 = gameLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_9 = gameLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_10 = gameLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_11 = gameLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_12 = gameLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_13 = gameLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_14 = gameLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_16 = gameLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_17 = gameLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_18 = gameLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_19 = gameLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_20 = gameLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_21 = gameLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_22 = gameLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_23 = gameLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_24 = gameLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_25 = gameLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_26 = gameLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_27 = gameLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_28 = gameLogic_io_spriteYPosition_28; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_29 = gameLogic_io_spriteYPosition_29; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_30 = gameLogic_io_spriteYPosition_30; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_31 = gameLogic_io_spriteYPosition_31; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_32 = gameLogic_io_spriteYPosition_32; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_33 = gameLogic_io_spriteYPosition_33; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_34 = gameLogic_io_spriteYPosition_34; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_35 = gameLogic_io_spriteYPosition_35; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_36 = gameLogic_io_spriteYPosition_36; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_37 = gameLogic_io_spriteYPosition_37; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_38 = gameLogic_io_spriteYPosition_38; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_39 = gameLogic_io_spriteYPosition_39; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_40 = gameLogic_io_spriteYPosition_40; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_41 = gameLogic_io_spriteYPosition_41; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_42 = gameLogic_io_spriteYPosition_42; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_43 = gameLogic_io_spriteYPosition_43; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_44 = gameLogic_io_spriteYPosition_44; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_45 = gameLogic_io_spriteYPosition_45; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_46 = gameLogic_io_spriteYPosition_46; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_47 = gameLogic_io_spriteYPosition_47; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_48 = gameLogic_io_spriteYPosition_48; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_49 = gameLogic_io_spriteYPosition_49; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_50 = gameLogic_io_spriteYPosition_50; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_51 = gameLogic_io_spriteYPosition_51; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_52 = gameLogic_io_spriteYPosition_52; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_53 = gameLogic_io_spriteYPosition_53; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_54 = gameLogic_io_spriteYPosition_54; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_55 = gameLogic_io_spriteYPosition_55; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_56 = gameLogic_io_spriteYPosition_56; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_57 = gameLogic_io_spriteYPosition_57; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_58 = gameLogic_io_spriteYPosition_58; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_59 = gameLogic_io_spriteYPosition_59; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_60 = gameLogic_io_spriteYPosition_60; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_61 = gameLogic_io_spriteYPosition_61; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_62 = gameLogic_io_spriteYPosition_62; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_63 = gameLogic_io_spriteYPosition_63; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteVisible_3 = gameLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_4 = gameLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_5 = gameLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_6 = gameLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_7 = gameLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_8 = gameLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_9 = gameLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_10 = gameLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_11 = gameLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_12 = gameLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_13 = gameLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_14 = gameLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_15 = gameLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_16 = gameLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_17 = gameLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_18 = gameLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_19 = gameLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_20 = gameLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_21 = gameLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_22 = gameLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_23 = gameLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_24 = gameLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_25 = gameLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_26 = gameLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_27 = gameLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_28 = gameLogic_io_spriteVisible_28; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_29 = gameLogic_io_spriteVisible_29; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_30 = gameLogic_io_spriteVisible_30; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_31 = gameLogic_io_spriteVisible_31; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_32 = gameLogic_io_spriteVisible_32; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_33 = gameLogic_io_spriteVisible_33; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_34 = gameLogic_io_spriteVisible_34; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_35 = gameLogic_io_spriteVisible_35; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_36 = gameLogic_io_spriteVisible_36; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_37 = gameLogic_io_spriteVisible_37; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_38 = gameLogic_io_spriteVisible_38; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_39 = gameLogic_io_spriteVisible_39; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_40 = gameLogic_io_spriteVisible_40; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_41 = gameLogic_io_spriteVisible_41; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_42 = gameLogic_io_spriteVisible_42; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_43 = gameLogic_io_spriteVisible_43; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_44 = gameLogic_io_spriteVisible_44; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_45 = gameLogic_io_spriteVisible_45; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_46 = gameLogic_io_spriteVisible_46; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_47 = gameLogic_io_spriteVisible_47; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_48 = gameLogic_io_spriteVisible_48; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_49 = gameLogic_io_spriteVisible_49; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_50 = gameLogic_io_spriteVisible_50; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_51 = gameLogic_io_spriteVisible_51; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_52 = gameLogic_io_spriteVisible_52; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_53 = gameLogic_io_spriteVisible_53; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_54 = gameLogic_io_spriteVisible_54; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_55 = gameLogic_io_spriteVisible_55; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_56 = gameLogic_io_spriteVisible_56; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_57 = gameLogic_io_spriteVisible_57; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_58 = gameLogic_io_spriteVisible_58; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_59 = gameLogic_io_spriteVisible_59; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_60 = gameLogic_io_spriteVisible_60; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_61 = gameLogic_io_spriteVisible_61; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_62 = gameLogic_io_spriteVisible_62; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_63 = gameLogic_io_spriteVisible_63; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_64 = gameLogic_io_spriteVisible_64; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_65 = gameLogic_io_spriteVisible_65; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_66 = gameLogic_io_spriteVisible_66; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_67 = gameLogic_io_spriteVisible_67; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_68 = gameLogic_io_spriteVisible_68; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_69 = gameLogic_io_spriteVisible_69; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_70 = gameLogic_io_spriteVisible_70; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_71 = gameLogic_io_spriteVisible_71; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_72 = gameLogic_io_spriteVisible_72; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_73 = gameLogic_io_spriteVisible_73; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_74 = gameLogic_io_spriteVisible_74; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_75 = gameLogic_io_spriteVisible_75; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_76 = gameLogic_io_spriteVisible_76; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_77 = gameLogic_io_spriteVisible_77; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_78 = gameLogic_io_spriteVisible_78; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_79 = gameLogic_io_spriteVisible_79; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_80 = gameLogic_io_spriteVisible_80; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_81 = gameLogic_io_spriteVisible_81; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_82 = gameLogic_io_spriteVisible_82; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_83 = gameLogic_io_spriteVisible_83; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_84 = gameLogic_io_spriteVisible_84; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_85 = gameLogic_io_spriteVisible_85; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_86 = gameLogic_io_spriteVisible_86; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_87 = gameLogic_io_spriteVisible_87; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_88 = gameLogic_io_spriteVisible_88; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_89 = gameLogic_io_spriteVisible_89; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_90 = gameLogic_io_spriteVisible_90; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_91 = gameLogic_io_spriteVisible_91; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_92 = gameLogic_io_spriteVisible_92; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_93 = gameLogic_io_spriteVisible_93; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_94 = gameLogic_io_spriteVisible_94; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_95 = gameLogic_io_spriteVisible_95; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_96 = gameLogic_io_spriteVisible_96; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_97 = gameLogic_io_spriteVisible_97; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_98 = gameLogic_io_spriteVisible_98; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_99 = gameLogic_io_spriteVisible_99; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_16 = gameLogic_io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_17 = gameLogic_io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_18 = gameLogic_io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_19 = gameLogic_io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_20 = gameLogic_io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_21 = gameLogic_io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_22 = gameLogic_io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_23 = gameLogic_io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_24 = gameLogic_io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_25 = gameLogic_io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_26 = gameLogic_io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_27 = gameLogic_io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_28 = gameLogic_io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_29 = gameLogic_io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_30 = gameLogic_io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_31 = gameLogic_io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_32 = gameLogic_io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_33 = gameLogic_io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_34 = gameLogic_io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_35 = gameLogic_io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_36 = gameLogic_io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_37 = gameLogic_io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_38 = gameLogic_io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_39 = gameLogic_io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_40 = gameLogic_io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_41 = gameLogic_io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_42 = gameLogic_io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_43 = gameLogic_io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_44 = gameLogic_io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_45 = gameLogic_io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_58 = gameLogic_io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_59 = gameLogic_io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_60 = gameLogic_io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpVertical_16 = gameLogic_io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_17 = gameLogic_io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_18 = gameLogic_io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_19 = gameLogic_io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_20 = gameLogic_io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_21 = gameLogic_io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_22 = gameLogic_io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_23 = gameLogic_io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_24 = gameLogic_io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_25 = gameLogic_io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_26 = gameLogic_io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_27 = gameLogic_io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_28 = gameLogic_io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_29 = gameLogic_io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_30 = gameLogic_io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_31 = gameLogic_io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_32 = gameLogic_io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_33 = gameLogic_io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_34 = gameLogic_io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_35 = gameLogic_io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_36 = gameLogic_io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_37 = gameLogic_io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_38 = gameLogic_io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_39 = gameLogic_io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_40 = gameLogic_io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_41 = gameLogic_io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_42 = gameLogic_io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_43 = gameLogic_io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_44 = gameLogic_io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_45 = gameLogic_io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_58 = gameLogic_io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_59 = gameLogic_io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_60 = gameLogic_io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_viewBoxX = gameLogic_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 138:32]
  assign graphicEngineVGA_io_viewBoxY = gameLogic_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 139:32]
  assign graphicEngineVGA_io_frameUpdateDone = gameLogic_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 148:39]
  assign soundEngine_clock = clock;
  assign soundEngine_reset = reset;
  assign gameLogic_clock = clock;
  assign gameLogic_reset = resetReleaseCounter == 22'h3d08ff ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameTop.scala 83:67 84:18 86:18]
  assign gameLogic_io_btnC = btnCState; // @[\\src\\main\\scala\\GameTop.scala 98:21]
  assign gameLogic_io_btnU = btnUState; // @[\\src\\main\\scala\\GameTop.scala 99:21]
  assign gameLogic_io_btnL = btnLState; // @[\\src\\main\\scala\\GameTop.scala 100:21]
  assign gameLogic_io_btnR = btnRState; // @[\\src\\main\\scala\\GameTop.scala 101:21]
  assign gameLogic_io_btnD = btnDState; // @[\\src\\main\\scala\\GameTop.scala 102:21]
  assign gameLogic_io_newFrame = graphicEngineVGA_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 147:25]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 68:32]
      debounceCounter <= 21'h0; // @[\\src\\main\\scala\\GameTop.scala 68:32]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 70:57]
      debounceCounter <= 21'h0; // @[\\src\\main\\scala\\GameTop.scala 71:21]
    end else begin
      debounceCounter <= _debounceCounter_T_1; // @[\\src\\main\\scala\\GameTop.scala 74:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 81:36]
      resetReleaseCounter <= 22'h0; // @[\\src\\main\\scala\\GameTop.scala 81:36]
    end else if (!(resetReleaseCounter == 22'h3d08ff)) begin // @[\\src\\main\\scala\\GameTop.scala 83:67]
      resetReleaseCounter <= _resetReleaseCounter_T_1; // @[\\src\\main\\scala\\GameTop.scala 87:25]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnCState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnCState_pipeReg_0 <= btnCState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnCState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnCState_pipeReg_1 <= btnCState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnCState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnCState_pipeReg_2 <= io_btnC; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 93:28]
      btnCState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 93:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 93:28]
      btnCState <= btnCState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 93:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_0 <= btnUState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_1 <= btnUState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_2 <= io_btnU; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 94:28]
      btnUState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 94:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 94:28]
      btnUState <= btnUState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 94:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_0 <= btnLState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_1 <= btnLState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_2 <= io_btnL; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 95:28]
      btnLState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 95:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 95:28]
      btnLState <= btnLState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 95:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_0 <= btnRState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_1 <= btnRState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_2 <= io_btnR; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 96:28]
      btnRState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 96:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 96:28]
      btnRState <= btnRState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 96:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_0 <= btnDState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_1 <= btnDState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_2 <= io_btnD; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 97:28]
      btnDState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 97:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 97:28]
      btnDState <= btnDState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 97:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounceCounter = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  resetReleaseCounter = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btnCState_pipeReg_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  btnCState_pipeReg_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  btnCState_pipeReg_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  btnCState = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  btnUState_pipeReg_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  btnUState_pipeReg_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  btnUState_pipeReg_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btnUState = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  btnLState_pipeReg_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  btnLState_pipeReg_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  btnLState_pipeReg_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btnLState = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  btnRState_pipeReg_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  btnRState_pipeReg_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  btnRState_pipeReg_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  btnRState = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  btnDState_pipeReg_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  btnDState_pipeReg_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  btnDState_pipeReg_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  btnDState = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input        clock,
  input        reset,
  input        io_btnC, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnU, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnL, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnR, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnD, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaRed, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaGreen, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaBlue, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_Hsync, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_Vsync, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_0, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_1, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_2, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_3, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_4, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_5, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_6, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_7, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_0, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_1, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_2, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_3, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_4, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_5, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_6, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_7, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_missingFrameError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_backBufferWriteError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_viewBoxOutOfRangeError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_soundOut // @[\\src\\main\\scala\\Top.scala 14:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  gameTop_clock; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_reset; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnC; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnU; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnL; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnR; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnD; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaRed; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaBlue; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaGreen; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_Hsync; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_Vsync; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_missingFrameError; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\Top.scala 44:23]
  reg  syncResetInput_REG; // @[\\src\\main\\scala\\Top.scala 49:48]
  reg  syncResetInput_REG_1; // @[\\src\\main\\scala\\Top.scala 49:40]
  reg  syncResetInput_REG_2; // @[\\src\\main\\scala\\Top.scala 49:32]
  reg  pipeResetReg_0; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_1; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_2; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_3; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_4; // @[\\src\\main\\scala\\Top.scala 54:25]
  wire [4:0] _gameTop_reset_T = {pipeResetReg_4,pipeResetReg_3,pipeResetReg_2,pipeResetReg_1,pipeResetReg_0}; // @[\\src\\main\\scala\\Top.scala 59:33]
  GameTop gameTop ( // @[\\src\\main\\scala\\Top.scala 44:23]
    .clock(gameTop_clock),
    .reset(gameTop_reset),
    .io_btnC(gameTop_io_btnC),
    .io_btnU(gameTop_io_btnU),
    .io_btnL(gameTop_io_btnL),
    .io_btnR(gameTop_io_btnR),
    .io_btnD(gameTop_io_btnD),
    .io_vgaRed(gameTop_io_vgaRed),
    .io_vgaBlue(gameTop_io_vgaBlue),
    .io_vgaGreen(gameTop_io_vgaGreen),
    .io_Hsync(gameTop_io_Hsync),
    .io_Vsync(gameTop_io_Vsync),
    .io_missingFrameError(gameTop_io_missingFrameError),
    .io_viewBoxOutOfRangeError(gameTop_io_viewBoxOutOfRangeError)
  );
  assign io_vgaRed = gameTop_io_vgaRed; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_vgaGreen = gameTop_io_vgaGreen; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_vgaBlue = gameTop_io_vgaBlue; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_Hsync = gameTop_io_Hsync; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_Vsync = gameTop_io_Vsync; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_0 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_1 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_2 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_3 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_4 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_5 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_6 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_7 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_missingFrameError = gameTop_io_missingFrameError; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_backBufferWriteError = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_viewBoxOutOfRangeError = gameTop_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_soundOut = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_clock = clock;
  assign gameTop_reset = |_gameTop_reset_T; // @[\\src\\main\\scala\\Top.scala 59:40]
  assign gameTop_io_btnC = io_btnC; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnU = io_btnU; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnL = io_btnL; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnR = io_btnR; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnD = io_btnD; // @[\\src\\main\\scala\\Top.scala 62:14]
  always @(posedge clock) begin
    syncResetInput_REG <= reset; // @[\\src\\main\\scala\\Top.scala 49:48]
    syncResetInput_REG_1 <= syncResetInput_REG; // @[\\src\\main\\scala\\Top.scala 49:40]
    syncResetInput_REG_2 <= syncResetInput_REG_1; // @[\\src\\main\\scala\\Top.scala 49:32]
    pipeResetReg_0 <= pipeResetReg_1; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_1 <= pipeResetReg_2; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_2 <= pipeResetReg_3; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_3 <= pipeResetReg_4; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_4 <= ~syncResetInput_REG_2; // @[\\src\\main\\scala\\Top.scala 49:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  syncResetInput_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  syncResetInput_REG_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  syncResetInput_REG_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pipeResetReg_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pipeResetReg_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pipeResetReg_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pipeResetReg_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pipeResetReg_4 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
