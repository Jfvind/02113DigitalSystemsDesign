module Memory(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_1(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_2(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_2.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_3(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_3.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_4(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_4.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_5(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_5.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_6(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_6.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_7(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_7.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_8(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_8.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_9(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_9.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_10(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_10.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_11(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_11.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_12(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_12.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_13(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_13.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_14(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_14.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_15(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_15.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_16(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_16.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_17(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_17.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_18(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_18.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_19(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_19.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_20(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_20.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_21(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_21.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_22(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_22.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_23(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_23.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_24(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_24.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_25(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_25.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_26(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_26.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_27(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_27.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_28(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_28.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_29(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_29.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_30(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_30.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_31(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_31.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_32(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_32.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_33(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_33.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_34(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_34.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_35(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_35.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_36(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_36.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_37(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_37.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_38(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_38.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_39(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_39.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_40(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_40.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_41(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_41.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_42(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_42.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_43(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_43.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_44(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_44.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_45(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_45.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_46(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_46.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_47(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_47.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_48(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_48.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_49(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_49.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_50(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_50.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_51(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_51.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_52(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_52.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_53(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_53.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_54(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_54.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_55(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_55.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_56(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_56.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_57(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_57.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_58(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_58.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_59(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_59.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_60(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_60.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_61(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_61.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_62(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_62.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_63(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_63.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_64(
  input         clock,
  input  [10:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [5:0]  io_dataRead, // @[\\src\\main\\scala\\Memory.scala 48:14]
  input         io_writeEnable, // @[\\src\\main\\scala\\Memory.scala 48:14]
  input  [5:0]  io_dataWrite // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [10:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [5:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [5:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 57:26]
  RamSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(6)) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 57:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 63:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 58:21]
  assign ramsSpWf_we = io_writeEnable; // @[\\src\\main\\scala\\Memory.scala 59:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 60:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 61:22]
  assign ramsSpWf_di = io_dataWrite; // @[\\src\\main\\scala\\Memory.scala 62:20]
endmodule
module Memory_66(
  input         clock,
  input  [10:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [5:0]  io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [10:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [5:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [5:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(6), .LOAD_FILE("memory_init/backbuffer_init.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 6'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_67(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_68(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_69(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_2.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_70(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_3.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_71(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_4.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_72(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_5.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_73(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_6.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_74(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_7.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_75(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_8.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_76(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_9.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_77(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_10.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_78(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_11.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_79(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_12.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_80(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_13.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_81(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_14.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_82(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_15.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_83(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_16.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_84(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_17.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_85(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_18.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_86(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_19.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_87(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_20.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_88(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_21.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_89(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_22.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_90(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_23.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_91(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_24.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_92(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_25.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_93(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_26.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_94(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_27.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_95(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_28.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_96(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_29.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_97(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_30.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_98(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_31.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_99(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_32.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_100(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_33.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_101(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_34.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_102(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_35.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_103(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_36.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_104(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_37.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_105(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_38.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_106(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_39.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_107(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_40.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_108(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_41.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_109(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_42.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_110(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_43.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_111(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_44.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_112(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_45.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_113(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_46.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_114(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_47.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_115(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_48.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_116(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_49.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_117(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_50.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_118(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_51.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_119(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_52.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_120(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_53.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_121(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_54.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_122(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_55.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_123(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_56.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_124(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_57.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_125(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_58.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_126(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_59.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_127(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_60.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_128(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_61.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_129(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_62.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_130(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_63.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module MultiHotPriortyReductionTree(
  input  [5:0] io_dataInput_0, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_1, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_2, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_3, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_4, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_5, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_6, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_7, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_8, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_9, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_10, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_11, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_12, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_13, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_14, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_15, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_16, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_17, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_18, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_19, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_20, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_21, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_22, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_23, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_24, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_25, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_26, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_27, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_28, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_29, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_30, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_31, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_32, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_33, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_34, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_35, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_36, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_37, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_38, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_39, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_40, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_41, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_42, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_43, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_44, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_45, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_46, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_47, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_48, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_49, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_50, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_51, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_52, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_53, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_54, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_55, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_56, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_57, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_58, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_59, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_60, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_61, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_62, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_63, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_0, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_1, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_2, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_3, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_4, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_5, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_6, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_7, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_8, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_9, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_10, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_11, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_12, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_13, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_14, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_15, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_16, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_17, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_18, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_19, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_20, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_21, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_22, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_23, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_24, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_25, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_26, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_27, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_28, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_29, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_30, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_31, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_32, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_33, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_34, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_35, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_36, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_37, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_38, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_39, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_40, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_41, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_42, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_43, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_44, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_45, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_46, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_47, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_48, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_49, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_50, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_51, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_52, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_53, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_54, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_55, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_56, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_57, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_58, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_59, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_60, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_61, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_62, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_63, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  output [5:0] io_dataOutput, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  output       io_selectOutput // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
);
  wire  selectNodeOutputs_31 = io_selectInput_0 | io_selectInput_1; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_32 = io_selectInput_2 | io_selectInput_3; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_15 = selectNodeOutputs_31 | selectNodeOutputs_32; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_33 = io_selectInput_4 | io_selectInput_5; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_34 = io_selectInput_6 | io_selectInput_7; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_16 = selectNodeOutputs_33 | selectNodeOutputs_34; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_7 = selectNodeOutputs_15 | selectNodeOutputs_16; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_35 = io_selectInput_8 | io_selectInput_9; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_36 = io_selectInput_10 | io_selectInput_11; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_17 = selectNodeOutputs_35 | selectNodeOutputs_36; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_37 = io_selectInput_12 | io_selectInput_13; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_38 = io_selectInput_14 | io_selectInput_15; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_18 = selectNodeOutputs_37 | selectNodeOutputs_38; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_8 = selectNodeOutputs_17 | selectNodeOutputs_18; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_3 = selectNodeOutputs_7 | selectNodeOutputs_8; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_39 = io_selectInput_16 | io_selectInput_17; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_40 = io_selectInput_18 | io_selectInput_19; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_19 = selectNodeOutputs_39 | selectNodeOutputs_40; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_41 = io_selectInput_20 | io_selectInput_21; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_42 = io_selectInput_22 | io_selectInput_23; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_20 = selectNodeOutputs_41 | selectNodeOutputs_42; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_9 = selectNodeOutputs_19 | selectNodeOutputs_20; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_43 = io_selectInput_24 | io_selectInput_25; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_44 = io_selectInput_26 | io_selectInput_27; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_21 = selectNodeOutputs_43 | selectNodeOutputs_44; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_45 = io_selectInput_28 | io_selectInput_29; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_46 = io_selectInput_30 | io_selectInput_31; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_22 = selectNodeOutputs_45 | selectNodeOutputs_46; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_10 = selectNodeOutputs_21 | selectNodeOutputs_22; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_4 = selectNodeOutputs_9 | selectNodeOutputs_10; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_1 = selectNodeOutputs_3 | selectNodeOutputs_4; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_31 = io_selectInput_0 ? io_dataInput_0 : io_dataInput_1; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_32 = io_selectInput_2 ? io_dataInput_2 : io_dataInput_3; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_15 = selectNodeOutputs_31 ? dataNodeOutputs_31 : dataNodeOutputs_32; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_33 = io_selectInput_4 ? io_dataInput_4 : io_dataInput_5; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_34 = io_selectInput_6 ? io_dataInput_6 : io_dataInput_7; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_16 = selectNodeOutputs_33 ? dataNodeOutputs_33 : dataNodeOutputs_34; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_7 = selectNodeOutputs_15 ? dataNodeOutputs_15 : dataNodeOutputs_16; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_35 = io_selectInput_8 ? io_dataInput_8 : io_dataInput_9; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_36 = io_selectInput_10 ? io_dataInput_10 : io_dataInput_11; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_17 = selectNodeOutputs_35 ? dataNodeOutputs_35 : dataNodeOutputs_36; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_37 = io_selectInput_12 ? io_dataInput_12 : io_dataInput_13; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_38 = io_selectInput_14 ? io_dataInput_14 : io_dataInput_15; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_18 = selectNodeOutputs_37 ? dataNodeOutputs_37 : dataNodeOutputs_38; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_8 = selectNodeOutputs_17 ? dataNodeOutputs_17 : dataNodeOutputs_18; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_3 = selectNodeOutputs_7 ? dataNodeOutputs_7 : dataNodeOutputs_8; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_39 = io_selectInput_16 ? io_dataInput_16 : io_dataInput_17; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_40 = io_selectInput_18 ? io_dataInput_18 : io_dataInput_19; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_19 = selectNodeOutputs_39 ? dataNodeOutputs_39 : dataNodeOutputs_40; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_41 = io_selectInput_20 ? io_dataInput_20 : io_dataInput_21; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_42 = io_selectInput_22 ? io_dataInput_22 : io_dataInput_23; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_20 = selectNodeOutputs_41 ? dataNodeOutputs_41 : dataNodeOutputs_42; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_9 = selectNodeOutputs_19 ? dataNodeOutputs_19 : dataNodeOutputs_20; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_43 = io_selectInput_24 ? io_dataInput_24 : io_dataInput_25; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_44 = io_selectInput_26 ? io_dataInput_26 : io_dataInput_27; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_21 = selectNodeOutputs_43 ? dataNodeOutputs_43 : dataNodeOutputs_44; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_45 = io_selectInput_28 ? io_dataInput_28 : io_dataInput_29; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_46 = io_selectInput_30 ? io_dataInput_30 : io_dataInput_31; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_22 = selectNodeOutputs_45 ? dataNodeOutputs_45 : dataNodeOutputs_46; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_10 = selectNodeOutputs_21 ? dataNodeOutputs_21 : dataNodeOutputs_22; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_4 = selectNodeOutputs_9 ? dataNodeOutputs_9 : dataNodeOutputs_10; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_1 = selectNodeOutputs_3 ? dataNodeOutputs_3 : dataNodeOutputs_4; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_47 = io_selectInput_32 | io_selectInput_33; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_48 = io_selectInput_34 | io_selectInput_35; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_23 = selectNodeOutputs_47 | selectNodeOutputs_48; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_49 = io_selectInput_36 | io_selectInput_37; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_50 = io_selectInput_38 | io_selectInput_39; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_24 = selectNodeOutputs_49 | selectNodeOutputs_50; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_11 = selectNodeOutputs_23 | selectNodeOutputs_24; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_51 = io_selectInput_40 | io_selectInput_41; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_52 = io_selectInput_42 | io_selectInput_43; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_25 = selectNodeOutputs_51 | selectNodeOutputs_52; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_53 = io_selectInput_44 | io_selectInput_45; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_54 = io_selectInput_46 | io_selectInput_47; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_26 = selectNodeOutputs_53 | selectNodeOutputs_54; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_12 = selectNodeOutputs_25 | selectNodeOutputs_26; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_5 = selectNodeOutputs_11 | selectNodeOutputs_12; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_47 = io_selectInput_32 ? io_dataInput_32 : io_dataInput_33; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_48 = io_selectInput_34 ? io_dataInput_34 : io_dataInput_35; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_23 = selectNodeOutputs_47 ? dataNodeOutputs_47 : dataNodeOutputs_48; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_49 = io_selectInput_36 ? io_dataInput_36 : io_dataInput_37; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_50 = io_selectInput_38 ? io_dataInput_38 : io_dataInput_39; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_24 = selectNodeOutputs_49 ? dataNodeOutputs_49 : dataNodeOutputs_50; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_11 = selectNodeOutputs_23 ? dataNodeOutputs_23 : dataNodeOutputs_24; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_51 = io_selectInput_40 ? io_dataInput_40 : io_dataInput_41; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_52 = io_selectInput_42 ? io_dataInput_42 : io_dataInput_43; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_25 = selectNodeOutputs_51 ? dataNodeOutputs_51 : dataNodeOutputs_52; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_53 = io_selectInput_44 ? io_dataInput_44 : io_dataInput_45; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_54 = io_selectInput_46 ? io_dataInput_46 : io_dataInput_47; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_26 = selectNodeOutputs_53 ? dataNodeOutputs_53 : dataNodeOutputs_54; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_12 = selectNodeOutputs_25 ? dataNodeOutputs_25 : dataNodeOutputs_26; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_5 = selectNodeOutputs_11 ? dataNodeOutputs_11 : dataNodeOutputs_12; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_55 = io_selectInput_48 | io_selectInput_49; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_56 = io_selectInput_50 | io_selectInput_51; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_27 = selectNodeOutputs_55 | selectNodeOutputs_56; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_57 = io_selectInput_52 | io_selectInput_53; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_58 = io_selectInput_54 | io_selectInput_55; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_28 = selectNodeOutputs_57 | selectNodeOutputs_58; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_13 = selectNodeOutputs_27 | selectNodeOutputs_28; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_55 = io_selectInput_48 ? io_dataInput_48 : io_dataInput_49; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_56 = io_selectInput_50 ? io_dataInput_50 : io_dataInput_51; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_27 = selectNodeOutputs_55 ? dataNodeOutputs_55 : dataNodeOutputs_56; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_57 = io_selectInput_52 ? io_dataInput_52 : io_dataInput_53; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_58 = io_selectInput_54 ? io_dataInput_54 : io_dataInput_55; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_28 = selectNodeOutputs_57 ? dataNodeOutputs_57 : dataNodeOutputs_58; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_13 = selectNodeOutputs_27 ? dataNodeOutputs_27 : dataNodeOutputs_28; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_59 = io_selectInput_56 | io_selectInput_57; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_60 = io_selectInput_58 | io_selectInput_59; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_29 = selectNodeOutputs_59 | selectNodeOutputs_60; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_59 = io_selectInput_56 ? io_dataInput_56 : io_dataInput_57; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_60 = io_selectInput_58 ? io_dataInput_58 : io_dataInput_59; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_29 = selectNodeOutputs_59 ? dataNodeOutputs_59 : dataNodeOutputs_60; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_61 = io_selectInput_60 | io_selectInput_61; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_61 = io_selectInput_60 ? io_dataInput_60 : io_dataInput_61; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_62 = io_selectInput_62 ? io_dataInput_62 : io_dataInput_63; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_30 = selectNodeOutputs_61 ? dataNodeOutputs_61 : dataNodeOutputs_62; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_14 = selectNodeOutputs_29 ? dataNodeOutputs_29 : dataNodeOutputs_30; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_6 = selectNodeOutputs_13 ? dataNodeOutputs_13 : dataNodeOutputs_14; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_2 = selectNodeOutputs_5 ? dataNodeOutputs_5 : dataNodeOutputs_6; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_62 = io_selectInput_62 | io_selectInput_63; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_30 = selectNodeOutputs_61 | selectNodeOutputs_62; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_14 = selectNodeOutputs_29 | selectNodeOutputs_30; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_6 = selectNodeOutputs_13 | selectNodeOutputs_14; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_2 = selectNodeOutputs_5 | selectNodeOutputs_6; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  assign io_dataOutput = selectNodeOutputs_1 ? dataNodeOutputs_1 : dataNodeOutputs_2; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  assign io_selectOutput = selectNodeOutputs_1 | selectNodeOutputs_2; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
endmodule
module GraphicEngineVGA(
  input         clock,
  input         reset,
  input  [10:0] io_spriteXPosition_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_46, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_47, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_48, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_49, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_50, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_51, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_52, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_53, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_54, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_55, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_56, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_57, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_61, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_62, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_63, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_46, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_47, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_48, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_49, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_50, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_51, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_52, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_53, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_54, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_55, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_56, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_57, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_61, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_62, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_63, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_4, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_5, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_6, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_15, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_46, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_47, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_48, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_49, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_50, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_51, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_52, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_53, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_54, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_55, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_56, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_57, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_61, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_62, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_63, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_viewBoxX, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [8:0]  io_viewBoxY, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_newFrame, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_frameUpdateDone, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_missingFrameError, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_viewBoxOutOfRangeError, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaRed, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaBlue, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaGreen, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_Hsync, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_Vsync // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
`endif // RANDOMIZE_REG_INIT
  wire  backTileMemories_0_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_0_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_1_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_1_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_2_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_2_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_3_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_3_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_4_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_4_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_5_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_5_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_6_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_6_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_7_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_7_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_8_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_8_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_9_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_9_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_10_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_10_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_11_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_11_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_12_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_12_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_13_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_13_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_14_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_14_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_15_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_15_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_16_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_16_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_17_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_17_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_18_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_18_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_19_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_19_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_20_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_20_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_21_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_21_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_22_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_22_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_23_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_23_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_24_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_24_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_25_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_25_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_26_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_26_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_27_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_27_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_28_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_28_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_29_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_29_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_30_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_30_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_31_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_31_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_32_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_32_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_32_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_33_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_33_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_33_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_34_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_34_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_34_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_35_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_35_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_35_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_36_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_36_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_36_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_37_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_37_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_37_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_38_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_38_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_38_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_39_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_39_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_39_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_40_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_40_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_40_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_41_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_41_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_41_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_42_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_42_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_42_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_43_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_43_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_43_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_44_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_44_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_44_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_45_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_45_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_45_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_46_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_46_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_46_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_47_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_47_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_47_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_48_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_48_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_48_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_49_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_49_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_49_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_50_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_50_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_50_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_51_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_51_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_51_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_52_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_52_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_52_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_53_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_53_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_53_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_54_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_54_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_54_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_55_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_55_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_55_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_56_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_56_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_56_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_57_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_57_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_57_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_58_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_58_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_58_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_59_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_59_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_59_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_60_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_60_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_60_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_61_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_61_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_61_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_62_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_62_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_62_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_63_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_63_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_63_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backBufferMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [10:0] backBufferMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [5:0] backBufferMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire  backBufferMemory_io_writeEnable; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [5:0] backBufferMemory_io_dataWrite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire  backBufferShadowMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [10:0] backBufferShadowMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [5:0] backBufferShadowMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire  backBufferShadowMemory_io_writeEnable; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [5:0] backBufferShadowMemory_io_dataWrite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire  backBufferRestoreMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire [10:0] backBufferRestoreMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire [5:0] backBufferRestoreMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire  spriteMemories_0_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_0_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_1_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_1_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_2_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_2_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_3_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_3_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_4_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_4_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_5_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_5_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_6_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_6_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_7_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_7_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_8_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_8_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_9_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_9_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_10_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_10_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_11_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_11_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_12_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_12_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_13_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_13_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_14_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_14_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_15_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_15_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_16_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_16_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_17_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_17_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_18_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_18_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_19_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_19_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_20_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_20_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_21_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_21_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_22_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_22_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_23_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_23_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_24_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_24_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_25_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_25_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_26_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_26_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_27_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_27_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_28_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_28_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_29_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_29_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_30_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_30_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_31_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_31_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_32_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_32_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_32_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_33_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_33_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_33_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_34_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_34_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_34_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_35_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_35_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_35_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_36_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_36_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_36_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_37_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_37_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_37_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_38_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_38_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_38_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_39_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_39_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_39_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_40_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_40_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_40_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_41_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_41_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_41_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_42_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_42_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_42_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_43_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_43_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_43_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_44_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_44_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_44_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_45_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_45_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_45_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_46_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_46_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_46_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_47_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_47_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_47_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_48_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_48_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_48_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_49_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_49_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_49_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_50_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_50_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_50_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_51_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_51_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_51_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_52_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_52_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_52_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_53_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_53_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_53_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_54_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_54_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_54_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_55_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_55_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_55_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_56_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_56_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_56_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_57_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_57_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_57_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_58_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_58_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_58_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_59_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_59_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_59_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_60_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_60_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_60_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_61_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_61_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_61_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_62_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_62_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_62_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_63_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_63_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_63_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  reg [1:0] ScaleCounterReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
  reg [9:0] CounterXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
  reg [9:0] CounterYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
  wire  _T_2 = CounterYReg == 10'h20c; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 78:26]
  wire [9:0] _CounterYReg_T_1 = CounterYReg + 10'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 82:38]
  wire [9:0] _GEN_0 = CounterYReg == 10'h20c ? 10'h0 : _CounterYReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 78:131 79:23 82:23]
  wire [9:0] _CounterXReg_T_1 = CounterXReg + 10'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 85:36]
  wire  _GEN_4 = CounterXReg == 10'h31f & _T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129 71:15]
  wire [1:0] _ScaleCounterReg_T_1 = ScaleCounterReg + 2'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 88:42]
  wire  _GEN_8 = ScaleCounterReg == 2'h3 & _GEN_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 71:15 74:52]
  reg [11:0] backMemoryRestoreCounter; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
  wire  restoreEnabled = backMemoryRestoreCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:33]
  wire  run = restoreEnabled ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:70 209:9 213:9]
  wire  Hsync = CounterXReg >= 10'h290 & CounterXReg < 10'h2f0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 92:79]
  wire  Vsync = CounterYReg >= 10'h1ea & CounterYReg < 10'h1ec; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 93:79]
  reg  io_Hsync_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg [20:0] frameClockCount; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
  wire [20:0] _frameClockCount_T_2 = frameClockCount + 21'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 105:92]
  wire  preDisplayArea = frameClockCount >= 21'h199a1b; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 106:40]
  reg [10:0] spriteXPositionReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [9:0] spriteYPositionReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg  spriteVisibleReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  wire  _GEN_141 = io_newFrame ? 1'h0 : spriteVisibleReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_142 = io_newFrame ? 1'h0 : spriteVisibleReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_143 = io_newFrame ? 1'h0 : spriteVisibleReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_144 = io_newFrame ? io_spriteVisible_3 : spriteVisibleReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_145 = io_newFrame ? io_spriteVisible_4 : spriteVisibleReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_146 = io_newFrame ? io_spriteVisible_5 : spriteVisibleReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_147 = io_newFrame ? io_spriteVisible_6 : spriteVisibleReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_148 = io_newFrame ? io_spriteVisible_7 : spriteVisibleReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_149 = io_newFrame ? io_spriteVisible_8 : spriteVisibleReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_150 = io_newFrame ? io_spriteVisible_9 : spriteVisibleReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_151 = io_newFrame ? io_spriteVisible_10 : spriteVisibleReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_152 = io_newFrame ? io_spriteVisible_11 : spriteVisibleReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_153 = io_newFrame ? io_spriteVisible_12 : spriteVisibleReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_154 = io_newFrame ? io_spriteVisible_13 : spriteVisibleReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_155 = io_newFrame ? io_spriteVisible_14 : spriteVisibleReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_156 = io_newFrame ? io_spriteVisible_15 : spriteVisibleReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_157 = io_newFrame ? io_spriteVisible_16 : spriteVisibleReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_158 = io_newFrame ? io_spriteVisible_17 : spriteVisibleReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_159 = io_newFrame ? io_spriteVisible_18 : spriteVisibleReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_160 = io_newFrame ? io_spriteVisible_19 : spriteVisibleReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_161 = io_newFrame ? io_spriteVisible_20 : spriteVisibleReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_162 = io_newFrame ? io_spriteVisible_21 : spriteVisibleReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_163 = io_newFrame ? io_spriteVisible_22 : spriteVisibleReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_164 = io_newFrame ? io_spriteVisible_23 : spriteVisibleReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_165 = io_newFrame ? io_spriteVisible_24 : spriteVisibleReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_166 = io_newFrame ? io_spriteVisible_25 : spriteVisibleReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_167 = io_newFrame ? io_spriteVisible_26 : spriteVisibleReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_168 = io_newFrame ? io_spriteVisible_27 : spriteVisibleReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_169 = io_newFrame ? io_spriteVisible_28 : spriteVisibleReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_170 = io_newFrame ? io_spriteVisible_29 : spriteVisibleReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_171 = io_newFrame ? io_spriteVisible_30 : spriteVisibleReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_172 = io_newFrame ? io_spriteVisible_31 : spriteVisibleReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_173 = io_newFrame ? io_spriteVisible_32 : spriteVisibleReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_174 = io_newFrame ? io_spriteVisible_33 : spriteVisibleReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_175 = io_newFrame ? io_spriteVisible_34 : spriteVisibleReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_176 = io_newFrame ? io_spriteVisible_35 : spriteVisibleReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_177 = io_newFrame ? io_spriteVisible_36 : spriteVisibleReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_178 = io_newFrame ? io_spriteVisible_37 : spriteVisibleReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_179 = io_newFrame ? io_spriteVisible_38 : spriteVisibleReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_180 = io_newFrame ? io_spriteVisible_39 : spriteVisibleReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_181 = io_newFrame ? io_spriteVisible_40 : spriteVisibleReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_182 = io_newFrame ? io_spriteVisible_41 : spriteVisibleReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_183 = io_newFrame ? io_spriteVisible_42 : spriteVisibleReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_184 = io_newFrame ? io_spriteVisible_43 : spriteVisibleReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_185 = io_newFrame ? io_spriteVisible_44 : spriteVisibleReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_186 = io_newFrame ? io_spriteVisible_45 : spriteVisibleReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_187 = io_newFrame ? io_spriteVisible_46 : spriteVisibleReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_188 = io_newFrame ? io_spriteVisible_47 : spriteVisibleReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_189 = io_newFrame ? io_spriteVisible_48 : spriteVisibleReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_190 = io_newFrame ? io_spriteVisible_49 : spriteVisibleReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_191 = io_newFrame ? io_spriteVisible_50 : spriteVisibleReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_192 = io_newFrame ? io_spriteVisible_51 : spriteVisibleReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_193 = io_newFrame ? io_spriteVisible_52 : spriteVisibleReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_194 = io_newFrame ? io_spriteVisible_53 : spriteVisibleReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_195 = io_newFrame ? io_spriteVisible_54 : spriteVisibleReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_196 = io_newFrame ? io_spriteVisible_55 : spriteVisibleReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_197 = io_newFrame ? io_spriteVisible_56 : spriteVisibleReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_198 = io_newFrame ? io_spriteVisible_57 : spriteVisibleReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_199 = io_newFrame ? io_spriteVisible_58 : spriteVisibleReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_200 = io_newFrame ? io_spriteVisible_59 : spriteVisibleReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_201 = io_newFrame ? io_spriteVisible_60 : spriteVisibleReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_202 = io_newFrame ? io_spriteVisible_61 : spriteVisibleReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_203 = io_newFrame ? io_spriteVisible_62 : spriteVisibleReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_204 = io_newFrame ? io_spriteVisible_63 : spriteVisibleReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  reg  spriteScaleUpHorizontalReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpVerticalReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg [9:0] viewBoxXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
  reg [8:0] viewBoxYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
  reg  missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
  reg  viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
  wire [9:0] viewBoxXClipped = viewBoxXReg >= 10'h280 ? 10'h280 : viewBoxXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 137:28]
  wire [8:0] viewBoxYClipped = viewBoxYReg >= 9'h1e0 ? 9'h1e0 : viewBoxYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 138:28]
  wire [10:0] pixelXBack = CounterXReg + viewBoxXClipped; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 139:27]
  wire [9:0] _GEN_1692 = {{1'd0}, viewBoxYClipped}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 140:27]
  wire [10:0] pixelYBack = CounterYReg + _GEN_1692; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 140:27]
  wire  _GEN_591 = viewBoxXReg > 10'h280 | viewBoxYReg > 9'h1e0 | viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 141:51 142:31 130:42]
  reg  newFrameStikyReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
  wire  _GEN_592 = io_newFrame | newFrameStikyReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 148:21 149:22 147:33]
  reg  REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:16]
  wire  _GEN_594 = newFrameStikyReg & io_newFrame | missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 154:41 155:26 128:37]
  wire [10:0] _backTileMemories_0_io_address_T_2 = 6'h20 * pixelYBack[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:75]
  wire [10:0] _GEN_1693 = {{6'd0}, pixelXBack[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:62]
  wire [11:0] _backTileMemories_0_io_address_T_3 = _GEN_1693 + _backTileMemories_0_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:62]
  reg [6:0] backTileMemoryDataRead_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [11:0] backMemoryCopyCounter; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
  wire  _T_7 = backMemoryCopyCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 187:32]
  wire [11:0] _backMemoryCopyCounter_T_1 = backMemoryCopyCounter + 12'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 188:54]
  wire  copyEnabled = preDisplayArea & _T_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23 198:17]
  reg  copyEnabledReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 200:31]
  wire [11:0] _backMemoryRestoreCounter_T_1 = backMemoryRestoreCounter + 12'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 206:58]
  reg [10:0] backBufferShadowMemory_io_address_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:67]
  wire [10:0] _backBufferShadowMemory_io_address_T_2 = copyEnabled ? backMemoryCopyCounter[10:0] : 11'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:105]
  reg  backBufferShadowMemory_io_writeEnable_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:71]
  reg [10:0] backBufferMemory_io_address_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:61]
  wire [11:0] _backBufferMemory_io_address_T_3 = 6'h28 * pixelYBack[10:5]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:130]
  wire [11:0] _GEN_1757 = {{6'd0}, pixelXBack[10:5]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:117]
  wire [12:0] _backBufferMemory_io_address_T_4 = _GEN_1757 + _backBufferMemory_io_address_T_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:117]
  wire [12:0] _backBufferMemory_io_address_T_5 = copyEnabledReg ? {{2'd0}, backBufferMemory_io_address_REG} :
    _backBufferMemory_io_address_T_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:37]
  reg [5:0] fullBackgroundColor_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:56]
  wire [6:0] _GEN_605 = 6'h1 == fullBackgroundColor_REG ? backTileMemoryDataRead_1_REG : backTileMemoryDataRead_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_606 = 6'h2 == fullBackgroundColor_REG ? backTileMemoryDataRead_2_REG : _GEN_605; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_607 = 6'h3 == fullBackgroundColor_REG ? backTileMemoryDataRead_3_REG : _GEN_606; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_608 = 6'h4 == fullBackgroundColor_REG ? backTileMemoryDataRead_4_REG : _GEN_607; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_609 = 6'h5 == fullBackgroundColor_REG ? backTileMemoryDataRead_5_REG : _GEN_608; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_610 = 6'h6 == fullBackgroundColor_REG ? backTileMemoryDataRead_6_REG : _GEN_609; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_611 = 6'h7 == fullBackgroundColor_REG ? backTileMemoryDataRead_7_REG : _GEN_610; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_612 = 6'h8 == fullBackgroundColor_REG ? backTileMemoryDataRead_8_REG : _GEN_611; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_613 = 6'h9 == fullBackgroundColor_REG ? backTileMemoryDataRead_9_REG : _GEN_612; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_614 = 6'ha == fullBackgroundColor_REG ? backTileMemoryDataRead_10_REG : _GEN_613; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_615 = 6'hb == fullBackgroundColor_REG ? backTileMemoryDataRead_11_REG : _GEN_614; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_616 = 6'hc == fullBackgroundColor_REG ? backTileMemoryDataRead_12_REG : _GEN_615; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_617 = 6'hd == fullBackgroundColor_REG ? backTileMemoryDataRead_13_REG : _GEN_616; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_618 = 6'he == fullBackgroundColor_REG ? backTileMemoryDataRead_14_REG : _GEN_617; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_619 = 6'hf == fullBackgroundColor_REG ? backTileMemoryDataRead_15_REG : _GEN_618; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_620 = 6'h10 == fullBackgroundColor_REG ? backTileMemoryDataRead_16_REG : _GEN_619; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_621 = 6'h11 == fullBackgroundColor_REG ? backTileMemoryDataRead_17_REG : _GEN_620; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_622 = 6'h12 == fullBackgroundColor_REG ? backTileMemoryDataRead_18_REG : _GEN_621; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_623 = 6'h13 == fullBackgroundColor_REG ? backTileMemoryDataRead_19_REG : _GEN_622; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_624 = 6'h14 == fullBackgroundColor_REG ? backTileMemoryDataRead_20_REG : _GEN_623; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_625 = 6'h15 == fullBackgroundColor_REG ? backTileMemoryDataRead_21_REG : _GEN_624; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_626 = 6'h16 == fullBackgroundColor_REG ? backTileMemoryDataRead_22_REG : _GEN_625; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_627 = 6'h17 == fullBackgroundColor_REG ? backTileMemoryDataRead_23_REG : _GEN_626; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_628 = 6'h18 == fullBackgroundColor_REG ? backTileMemoryDataRead_24_REG : _GEN_627; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_629 = 6'h19 == fullBackgroundColor_REG ? backTileMemoryDataRead_25_REG : _GEN_628; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_630 = 6'h1a == fullBackgroundColor_REG ? backTileMemoryDataRead_26_REG : _GEN_629; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_631 = 6'h1b == fullBackgroundColor_REG ? backTileMemoryDataRead_27_REG : _GEN_630; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_632 = 6'h1c == fullBackgroundColor_REG ? backTileMemoryDataRead_28_REG : _GEN_631; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_633 = 6'h1d == fullBackgroundColor_REG ? backTileMemoryDataRead_29_REG : _GEN_632; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_634 = 6'h1e == fullBackgroundColor_REG ? backTileMemoryDataRead_30_REG : _GEN_633; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_635 = 6'h1f == fullBackgroundColor_REG ? backTileMemoryDataRead_31_REG : _GEN_634; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_636 = 6'h20 == fullBackgroundColor_REG ? backTileMemoryDataRead_32_REG : _GEN_635; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_637 = 6'h21 == fullBackgroundColor_REG ? backTileMemoryDataRead_33_REG : _GEN_636; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_638 = 6'h22 == fullBackgroundColor_REG ? backTileMemoryDataRead_34_REG : _GEN_637; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_639 = 6'h23 == fullBackgroundColor_REG ? backTileMemoryDataRead_35_REG : _GEN_638; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_640 = 6'h24 == fullBackgroundColor_REG ? backTileMemoryDataRead_36_REG : _GEN_639; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_641 = 6'h25 == fullBackgroundColor_REG ? backTileMemoryDataRead_37_REG : _GEN_640; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_642 = 6'h26 == fullBackgroundColor_REG ? backTileMemoryDataRead_38_REG : _GEN_641; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_643 = 6'h27 == fullBackgroundColor_REG ? backTileMemoryDataRead_39_REG : _GEN_642; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_644 = 6'h28 == fullBackgroundColor_REG ? backTileMemoryDataRead_40_REG : _GEN_643; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_645 = 6'h29 == fullBackgroundColor_REG ? backTileMemoryDataRead_41_REG : _GEN_644; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_646 = 6'h2a == fullBackgroundColor_REG ? backTileMemoryDataRead_42_REG : _GEN_645; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_647 = 6'h2b == fullBackgroundColor_REG ? backTileMemoryDataRead_43_REG : _GEN_646; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_648 = 6'h2c == fullBackgroundColor_REG ? backTileMemoryDataRead_44_REG : _GEN_647; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_649 = 6'h2d == fullBackgroundColor_REG ? backTileMemoryDataRead_45_REG : _GEN_648; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_650 = 6'h2e == fullBackgroundColor_REG ? backTileMemoryDataRead_46_REG : _GEN_649; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_651 = 6'h2f == fullBackgroundColor_REG ? backTileMemoryDataRead_47_REG : _GEN_650; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_652 = 6'h30 == fullBackgroundColor_REG ? backTileMemoryDataRead_48_REG : _GEN_651; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_653 = 6'h31 == fullBackgroundColor_REG ? backTileMemoryDataRead_49_REG : _GEN_652; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_654 = 6'h32 == fullBackgroundColor_REG ? backTileMemoryDataRead_50_REG : _GEN_653; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_655 = 6'h33 == fullBackgroundColor_REG ? backTileMemoryDataRead_51_REG : _GEN_654; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_656 = 6'h34 == fullBackgroundColor_REG ? backTileMemoryDataRead_52_REG : _GEN_655; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_657 = 6'h35 == fullBackgroundColor_REG ? backTileMemoryDataRead_53_REG : _GEN_656; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_658 = 6'h36 == fullBackgroundColor_REG ? backTileMemoryDataRead_54_REG : _GEN_657; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_659 = 6'h37 == fullBackgroundColor_REG ? backTileMemoryDataRead_55_REG : _GEN_658; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_660 = 6'h38 == fullBackgroundColor_REG ? backTileMemoryDataRead_56_REG : _GEN_659; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_661 = 6'h39 == fullBackgroundColor_REG ? backTileMemoryDataRead_57_REG : _GEN_660; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_662 = 6'h3a == fullBackgroundColor_REG ? backTileMemoryDataRead_58_REG : _GEN_661; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_663 = 6'h3b == fullBackgroundColor_REG ? backTileMemoryDataRead_59_REG : _GEN_662; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_664 = 6'h3c == fullBackgroundColor_REG ? backTileMemoryDataRead_60_REG : _GEN_663; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_665 = 6'h3d == fullBackgroundColor_REG ? backTileMemoryDataRead_61_REG : _GEN_664; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_666 = 6'h3e == fullBackgroundColor_REG ? backTileMemoryDataRead_62_REG : _GEN_665; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] fullBackgroundColor = 6'h3f == fullBackgroundColor_REG ? backTileMemoryDataRead_63_REG : _GEN_666; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  reg [5:0] pixelColorBack; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 245:31]
  wire [10:0] _inSpriteXValue_T_1 = {1'h0,CounterXReg}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:47]
  wire [11:0] inSpriteXValue = $signed(_inSpriteXValue_T_1) - 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_0 = $signed(inSpriteXValue) >= 12'sh0 & $signed(inSpriteXValue) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_674 = {{1{inSpriteXValue[11]}},inSpriteXValue}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _inSpriteYValue_T_1 = {1'h0,CounterYReg}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:47]
  wire [11:0] inSpriteYValue = $signed(_inSpriteYValue_T_1) - 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_0 = inSpriteYValue[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_0 = $signed(inSpriteYPreScaled_0) >= 11'sh0 & $signed(inSpriteYPreScaled_0) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_682 = {{1{inSpriteYPreScaled_0[10]}},inSpriteYPreScaled_0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_3 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_3); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_3 = $signed(inSpriteXValue_3) >= 12'sh0 & $signed(inSpriteXValue_3) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_722 = {{1{inSpriteXValue_3[11]}},inSpriteXValue_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1761 = {{1{spriteYPositionReg_3[9]}},spriteYPositionReg_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_3 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1761); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_3 = inSpriteYValue_3[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_3 = $signed(inSpriteYPreScaled_3) >= 11'sh0 & $signed(inSpriteYPreScaled_3) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_730 = {{1{inSpriteYPreScaled_3[10]}},inSpriteYPreScaled_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_7 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_7); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_7 = $signed(inSpriteXValue_7) >= 12'sh0 & $signed(inSpriteXValue_7) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_786 = {{1{inSpriteXValue_7[11]}},inSpriteXValue_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1766 = {{1{spriteYPositionReg_7[9]}},spriteYPositionReg_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_7 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1766); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_7 = inSpriteYValue_7[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_7 = $signed(inSpriteYPreScaled_7) >= 11'sh0 & $signed(inSpriteYPreScaled_7) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_794 = {{1{inSpriteYPreScaled_7[10]}},inSpriteYPreScaled_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_8 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_8); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_8 = $signed(inSpriteXValue_8) >= 12'sh0 & $signed(inSpriteXValue_8) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_802 = {{1{inSpriteXValue_8[11]}},inSpriteXValue_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1768 = {{1{spriteYPositionReg_8[9]}},spriteYPositionReg_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_8 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1768); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_8 = inSpriteYValue_8[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_8 = $signed(inSpriteYPreScaled_8) >= 11'sh0 & $signed(inSpriteYPreScaled_8) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_810 = {{1{inSpriteYPreScaled_8[10]}},inSpriteYPreScaled_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_9 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_9); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_9 = $signed(inSpriteXValue_9) >= 12'sh0 & $signed(inSpriteXValue_9) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_818 = {{1{inSpriteXValue_9[11]}},inSpriteXValue_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1770 = {{1{spriteYPositionReg_9[9]}},spriteYPositionReg_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_9 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1770); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_9 = inSpriteYValue_9[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_9 = $signed(inSpriteYPreScaled_9) >= 11'sh0 & $signed(inSpriteYPreScaled_9) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_826 = {{1{inSpriteYPreScaled_9[10]}},inSpriteYPreScaled_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_10 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_10); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_10 = $signed(inSpriteXValue_10) >= 12'sh0 & $signed(inSpriteXValue_10) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_834 = {{1{inSpriteXValue_10[11]}},inSpriteXValue_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1772 = {{1{spriteYPositionReg_10[9]}},spriteYPositionReg_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_10 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1772); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_10 = inSpriteYValue_10[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_10 = $signed(inSpriteYPreScaled_10) >= 11'sh0 & $signed(inSpriteYPreScaled_10) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_842 = {{1{inSpriteYPreScaled_10[10]}},inSpriteYPreScaled_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_11 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_11); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_11 = $signed(inSpriteXValue_11) >= 12'sh0 & $signed(inSpriteXValue_11) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_850 = {{1{inSpriteXValue_11[11]}},inSpriteXValue_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1774 = {{1{spriteYPositionReg_11[9]}},spriteYPositionReg_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_11 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1774); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_11 = inSpriteYValue_11[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_11 = $signed(inSpriteYPreScaled_11) >= 11'sh0 & $signed(inSpriteYPreScaled_11) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_858 = {{1{inSpriteYPreScaled_11[10]}},inSpriteYPreScaled_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_12 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_12); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_12 = $signed(inSpriteXValue_12) >= 12'sh0 & $signed(inSpriteXValue_12) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_866 = {{1{inSpriteXValue_12[11]}},inSpriteXValue_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1776 = {{1{spriteYPositionReg_12[9]}},spriteYPositionReg_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_12 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1776); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_12 = inSpriteYValue_12[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_12 = $signed(inSpriteYPreScaled_12) >= 11'sh0 & $signed(inSpriteYPreScaled_12) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_874 = {{1{inSpriteYPreScaled_12[10]}},inSpriteYPreScaled_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_13 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_13); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_13 = $signed(inSpriteXValue_13) >= 12'sh0 & $signed(inSpriteXValue_13) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_882 = {{1{inSpriteXValue_13[11]}},inSpriteXValue_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1778 = {{1{spriteYPositionReg_13[9]}},spriteYPositionReg_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_13 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1778); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_13 = inSpriteYValue_13[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_13 = $signed(inSpriteYPreScaled_13) >= 11'sh0 & $signed(inSpriteYPreScaled_13) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_890 = {{1{inSpriteYPreScaled_13[10]}},inSpriteYPreScaled_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_14 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_14); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_14 = $signed(inSpriteXValue_14) >= 12'sh0 & $signed(inSpriteXValue_14) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_898 = {{1{inSpriteXValue_14[11]}},inSpriteXValue_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1780 = {{1{spriteYPositionReg_14[9]}},spriteYPositionReg_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_14 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1780); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_14 = inSpriteYValue_14[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_14 = $signed(inSpriteYPreScaled_14) >= 11'sh0 & $signed(inSpriteYPreScaled_14) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_906 = {{1{inSpriteYPreScaled_14[10]}},inSpriteYPreScaled_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_16 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_16); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_16_T = $signed(inSpriteXValue_16) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_16_T_4 = inSpriteXValue_16[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_16_T_8 = _inSpriteHorizontal_16_T & $signed(inSpriteXValue_16) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_16_T_5 = {$signed(inSpriteXValue_16), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_16_T_14 = _inSpriteHorizontal_16_T & $signed(inSpriteXValue_16) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_928 = spriteScaleUpHorizontalReg_16 ? $signed({{2{_inSpriteX_16_T_4[10]}},_inSpriteX_16_T_4}) :
    $signed(_inSpriteX_16_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_929 = spriteScaleUpHorizontalReg_16 ? _inSpriteHorizontal_16_T_8 : _inSpriteHorizontal_16_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_930 = ~spriteScaleUpHorizontalReg_16 ? $signed({{1{inSpriteXValue_16[11]}},inSpriteXValue_16}) :
    $signed(_GEN_928); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_16 = ~spriteScaleUpHorizontalReg_16 ? $signed(inSpriteXValue_16) >= 12'sh0 & $signed(
    inSpriteXValue_16) < 12'sh20 : _GEN_929; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1783 = {{1{spriteYPositionReg_16[9]}},spriteYPositionReg_16}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_16 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1783); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_16 = inSpriteYValue_16[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_16_T = $signed(inSpriteYPreScaled_16) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_16_T_4 = inSpriteYPreScaled_16[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_16_T_8 = _inSpriteVertical_16_T & $signed(inSpriteYPreScaled_16) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_16_T_5 = {$signed(inSpriteYPreScaled_16), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_16_T_14 = _inSpriteVertical_16_T & $signed(inSpriteYPreScaled_16) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_936 = spriteScaleUpVerticalReg_16 ? $signed({{2{_inSpriteY_16_T_4[9]}},_inSpriteY_16_T_4}) : $signed(
    _inSpriteY_16_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_937 = spriteScaleUpVerticalReg_16 ? _inSpriteVertical_16_T_8 : _inSpriteVertical_16_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_938 = ~spriteScaleUpVerticalReg_16 ? $signed({{1{inSpriteYPreScaled_16[10]}},inSpriteYPreScaled_16})
     : $signed(_GEN_936); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_16 = ~spriteScaleUpVerticalReg_16 ? $signed(inSpriteYPreScaled_16) >= 11'sh0 & $signed(
    inSpriteYPreScaled_16) < 11'sh20 : _GEN_937; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_17 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_17); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_17_T = $signed(inSpriteXValue_17) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_17_T_4 = inSpriteXValue_17[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_17_T_8 = _inSpriteHorizontal_17_T & $signed(inSpriteXValue_17) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_17_T_5 = {$signed(inSpriteXValue_17), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_17_T_14 = _inSpriteHorizontal_17_T & $signed(inSpriteXValue_17) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_944 = spriteScaleUpHorizontalReg_17 ? $signed({{2{_inSpriteX_17_T_4[10]}},_inSpriteX_17_T_4}) :
    $signed(_inSpriteX_17_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_945 = spriteScaleUpHorizontalReg_17 ? _inSpriteHorizontal_17_T_8 : _inSpriteHorizontal_17_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_946 = ~spriteScaleUpHorizontalReg_17 ? $signed({{1{inSpriteXValue_17[11]}},inSpriteXValue_17}) :
    $signed(_GEN_944); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_17 = ~spriteScaleUpHorizontalReg_17 ? $signed(inSpriteXValue_17) >= 12'sh0 & $signed(
    inSpriteXValue_17) < 12'sh20 : _GEN_945; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1785 = {{1{spriteYPositionReg_17[9]}},spriteYPositionReg_17}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_17 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1785); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_17 = inSpriteYValue_17[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_17_T = $signed(inSpriteYPreScaled_17) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_17_T_4 = inSpriteYPreScaled_17[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_17_T_8 = _inSpriteVertical_17_T & $signed(inSpriteYPreScaled_17) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_17_T_5 = {$signed(inSpriteYPreScaled_17), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_17_T_14 = _inSpriteVertical_17_T & $signed(inSpriteYPreScaled_17) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_952 = spriteScaleUpVerticalReg_17 ? $signed({{2{_inSpriteY_17_T_4[9]}},_inSpriteY_17_T_4}) : $signed(
    _inSpriteY_17_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_953 = spriteScaleUpVerticalReg_17 ? _inSpriteVertical_17_T_8 : _inSpriteVertical_17_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_954 = ~spriteScaleUpVerticalReg_17 ? $signed({{1{inSpriteYPreScaled_17[10]}},inSpriteYPreScaled_17})
     : $signed(_GEN_952); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_17 = ~spriteScaleUpVerticalReg_17 ? $signed(inSpriteYPreScaled_17) >= 11'sh0 & $signed(
    inSpriteYPreScaled_17) < 11'sh20 : _GEN_953; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_18 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_18); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_18_T = $signed(inSpriteXValue_18) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_18_T_4 = inSpriteXValue_18[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_18_T_8 = _inSpriteHorizontal_18_T & $signed(inSpriteXValue_18) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_18_T_5 = {$signed(inSpriteXValue_18), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_18_T_14 = _inSpriteHorizontal_18_T & $signed(inSpriteXValue_18) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_960 = spriteScaleUpHorizontalReg_18 ? $signed({{2{_inSpriteX_18_T_4[10]}},_inSpriteX_18_T_4}) :
    $signed(_inSpriteX_18_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_961 = spriteScaleUpHorizontalReg_18 ? _inSpriteHorizontal_18_T_8 : _inSpriteHorizontal_18_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_962 = ~spriteScaleUpHorizontalReg_18 ? $signed({{1{inSpriteXValue_18[11]}},inSpriteXValue_18}) :
    $signed(_GEN_960); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_18 = ~spriteScaleUpHorizontalReg_18 ? $signed(inSpriteXValue_18) >= 12'sh0 & $signed(
    inSpriteXValue_18) < 12'sh20 : _GEN_961; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1787 = {{1{spriteYPositionReg_18[9]}},spriteYPositionReg_18}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_18 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1787); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_18 = inSpriteYValue_18[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_18_T = $signed(inSpriteYPreScaled_18) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_18_T_4 = inSpriteYPreScaled_18[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_18_T_8 = _inSpriteVertical_18_T & $signed(inSpriteYPreScaled_18) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_18_T_5 = {$signed(inSpriteYPreScaled_18), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_18_T_14 = _inSpriteVertical_18_T & $signed(inSpriteYPreScaled_18) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_968 = spriteScaleUpVerticalReg_18 ? $signed({{2{_inSpriteY_18_T_4[9]}},_inSpriteY_18_T_4}) : $signed(
    _inSpriteY_18_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_969 = spriteScaleUpVerticalReg_18 ? _inSpriteVertical_18_T_8 : _inSpriteVertical_18_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_970 = ~spriteScaleUpVerticalReg_18 ? $signed({{1{inSpriteYPreScaled_18[10]}},inSpriteYPreScaled_18})
     : $signed(_GEN_968); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_18 = ~spriteScaleUpVerticalReg_18 ? $signed(inSpriteYPreScaled_18) >= 11'sh0 & $signed(
    inSpriteYPreScaled_18) < 11'sh20 : _GEN_969; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_19 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_19); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_19_T = $signed(inSpriteXValue_19) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_19_T_4 = inSpriteXValue_19[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_19_T_8 = _inSpriteHorizontal_19_T & $signed(inSpriteXValue_19) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_19_T_5 = {$signed(inSpriteXValue_19), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_19_T_14 = _inSpriteHorizontal_19_T & $signed(inSpriteXValue_19) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_976 = spriteScaleUpHorizontalReg_19 ? $signed({{2{_inSpriteX_19_T_4[10]}},_inSpriteX_19_T_4}) :
    $signed(_inSpriteX_19_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_977 = spriteScaleUpHorizontalReg_19 ? _inSpriteHorizontal_19_T_8 : _inSpriteHorizontal_19_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_978 = ~spriteScaleUpHorizontalReg_19 ? $signed({{1{inSpriteXValue_19[11]}},inSpriteXValue_19}) :
    $signed(_GEN_976); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_19 = ~spriteScaleUpHorizontalReg_19 ? $signed(inSpriteXValue_19) >= 12'sh0 & $signed(
    inSpriteXValue_19) < 12'sh20 : _GEN_977; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1789 = {{1{spriteYPositionReg_19[9]}},spriteYPositionReg_19}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_19 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1789); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_19 = inSpriteYValue_19[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_19_T = $signed(inSpriteYPreScaled_19) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_19_T_4 = inSpriteYPreScaled_19[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_19_T_8 = _inSpriteVertical_19_T & $signed(inSpriteYPreScaled_19) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_19_T_5 = {$signed(inSpriteYPreScaled_19), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_19_T_14 = _inSpriteVertical_19_T & $signed(inSpriteYPreScaled_19) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_984 = spriteScaleUpVerticalReg_19 ? $signed({{2{_inSpriteY_19_T_4[9]}},_inSpriteY_19_T_4}) : $signed(
    _inSpriteY_19_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_985 = spriteScaleUpVerticalReg_19 ? _inSpriteVertical_19_T_8 : _inSpriteVertical_19_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_986 = ~spriteScaleUpVerticalReg_19 ? $signed({{1{inSpriteYPreScaled_19[10]}},inSpriteYPreScaled_19})
     : $signed(_GEN_984); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_19 = ~spriteScaleUpVerticalReg_19 ? $signed(inSpriteYPreScaled_19) >= 11'sh0 & $signed(
    inSpriteYPreScaled_19) < 11'sh20 : _GEN_985; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_20 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_20); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_20_T = $signed(inSpriteXValue_20) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_20_T_4 = inSpriteXValue_20[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_20_T_8 = _inSpriteHorizontal_20_T & $signed(inSpriteXValue_20) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_20_T_5 = {$signed(inSpriteXValue_20), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_20_T_14 = _inSpriteHorizontal_20_T & $signed(inSpriteXValue_20) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_992 = spriteScaleUpHorizontalReg_20 ? $signed({{2{_inSpriteX_20_T_4[10]}},_inSpriteX_20_T_4}) :
    $signed(_inSpriteX_20_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_993 = spriteScaleUpHorizontalReg_20 ? _inSpriteHorizontal_20_T_8 : _inSpriteHorizontal_20_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_994 = ~spriteScaleUpHorizontalReg_20 ? $signed({{1{inSpriteXValue_20[11]}},inSpriteXValue_20}) :
    $signed(_GEN_992); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_20 = ~spriteScaleUpHorizontalReg_20 ? $signed(inSpriteXValue_20) >= 12'sh0 & $signed(
    inSpriteXValue_20) < 12'sh20 : _GEN_993; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1791 = {{1{spriteYPositionReg_20[9]}},spriteYPositionReg_20}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_20 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1791); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_20 = inSpriteYValue_20[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_20_T = $signed(inSpriteYPreScaled_20) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_20_T_4 = inSpriteYPreScaled_20[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_20_T_8 = _inSpriteVertical_20_T & $signed(inSpriteYPreScaled_20) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_20_T_5 = {$signed(inSpriteYPreScaled_20), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_20_T_14 = _inSpriteVertical_20_T & $signed(inSpriteYPreScaled_20) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1000 = spriteScaleUpVerticalReg_20 ? $signed({{2{_inSpriteY_20_T_4[9]}},_inSpriteY_20_T_4}) :
    $signed(_inSpriteY_20_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1001 = spriteScaleUpVerticalReg_20 ? _inSpriteVertical_20_T_8 : _inSpriteVertical_20_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1002 = ~spriteScaleUpVerticalReg_20 ? $signed({{1{inSpriteYPreScaled_20[10]}},inSpriteYPreScaled_20})
     : $signed(_GEN_1000); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_20 = ~spriteScaleUpVerticalReg_20 ? $signed(inSpriteYPreScaled_20) >= 11'sh0 & $signed(
    inSpriteYPreScaled_20) < 11'sh20 : _GEN_1001; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_21 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_21); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_21_T = $signed(inSpriteXValue_21) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_21_T_4 = inSpriteXValue_21[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_21_T_8 = _inSpriteHorizontal_21_T & $signed(inSpriteXValue_21) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_21_T_5 = {$signed(inSpriteXValue_21), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_21_T_14 = _inSpriteHorizontal_21_T & $signed(inSpriteXValue_21) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1008 = spriteScaleUpHorizontalReg_21 ? $signed({{2{_inSpriteX_21_T_4[10]}},_inSpriteX_21_T_4}) :
    $signed(_inSpriteX_21_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1009 = spriteScaleUpHorizontalReg_21 ? _inSpriteHorizontal_21_T_8 : _inSpriteHorizontal_21_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1010 = ~spriteScaleUpHorizontalReg_21 ? $signed({{1{inSpriteXValue_21[11]}},inSpriteXValue_21}) :
    $signed(_GEN_1008); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_21 = ~spriteScaleUpHorizontalReg_21 ? $signed(inSpriteXValue_21) >= 12'sh0 & $signed(
    inSpriteXValue_21) < 12'sh20 : _GEN_1009; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1793 = {{1{spriteYPositionReg_21[9]}},spriteYPositionReg_21}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_21 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1793); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_21 = inSpriteYValue_21[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_21_T = $signed(inSpriteYPreScaled_21) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_21_T_4 = inSpriteYPreScaled_21[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_21_T_8 = _inSpriteVertical_21_T & $signed(inSpriteYPreScaled_21) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_21_T_5 = {$signed(inSpriteYPreScaled_21), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_21_T_14 = _inSpriteVertical_21_T & $signed(inSpriteYPreScaled_21) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1016 = spriteScaleUpVerticalReg_21 ? $signed({{2{_inSpriteY_21_T_4[9]}},_inSpriteY_21_T_4}) :
    $signed(_inSpriteY_21_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1017 = spriteScaleUpVerticalReg_21 ? _inSpriteVertical_21_T_8 : _inSpriteVertical_21_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1018 = ~spriteScaleUpVerticalReg_21 ? $signed({{1{inSpriteYPreScaled_21[10]}},inSpriteYPreScaled_21})
     : $signed(_GEN_1016); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_21 = ~spriteScaleUpVerticalReg_21 ? $signed(inSpriteYPreScaled_21) >= 11'sh0 & $signed(
    inSpriteYPreScaled_21) < 11'sh20 : _GEN_1017; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_22 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_22); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_22_T = $signed(inSpriteXValue_22) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_22_T_4 = inSpriteXValue_22[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_22_T_8 = _inSpriteHorizontal_22_T & $signed(inSpriteXValue_22) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_22_T_5 = {$signed(inSpriteXValue_22), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_22_T_14 = _inSpriteHorizontal_22_T & $signed(inSpriteXValue_22) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1024 = spriteScaleUpHorizontalReg_22 ? $signed({{2{_inSpriteX_22_T_4[10]}},_inSpriteX_22_T_4}) :
    $signed(_inSpriteX_22_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1025 = spriteScaleUpHorizontalReg_22 ? _inSpriteHorizontal_22_T_8 : _inSpriteHorizontal_22_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1026 = ~spriteScaleUpHorizontalReg_22 ? $signed({{1{inSpriteXValue_22[11]}},inSpriteXValue_22}) :
    $signed(_GEN_1024); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_22 = ~spriteScaleUpHorizontalReg_22 ? $signed(inSpriteXValue_22) >= 12'sh0 & $signed(
    inSpriteXValue_22) < 12'sh20 : _GEN_1025; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1795 = {{1{spriteYPositionReg_22[9]}},spriteYPositionReg_22}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_22 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1795); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_22 = inSpriteYValue_22[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_22_T = $signed(inSpriteYPreScaled_22) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_22_T_4 = inSpriteYPreScaled_22[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_22_T_8 = _inSpriteVertical_22_T & $signed(inSpriteYPreScaled_22) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_22_T_5 = {$signed(inSpriteYPreScaled_22), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_22_T_14 = _inSpriteVertical_22_T & $signed(inSpriteYPreScaled_22) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1032 = spriteScaleUpVerticalReg_22 ? $signed({{2{_inSpriteY_22_T_4[9]}},_inSpriteY_22_T_4}) :
    $signed(_inSpriteY_22_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1033 = spriteScaleUpVerticalReg_22 ? _inSpriteVertical_22_T_8 : _inSpriteVertical_22_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1034 = ~spriteScaleUpVerticalReg_22 ? $signed({{1{inSpriteYPreScaled_22[10]}},inSpriteYPreScaled_22})
     : $signed(_GEN_1032); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_22 = ~spriteScaleUpVerticalReg_22 ? $signed(inSpriteYPreScaled_22) >= 11'sh0 & $signed(
    inSpriteYPreScaled_22) < 11'sh20 : _GEN_1033; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_23 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_23); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_23_T = $signed(inSpriteXValue_23) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_23_T_4 = inSpriteXValue_23[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_23_T_8 = _inSpriteHorizontal_23_T & $signed(inSpriteXValue_23) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_23_T_5 = {$signed(inSpriteXValue_23), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_23_T_14 = _inSpriteHorizontal_23_T & $signed(inSpriteXValue_23) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1040 = spriteScaleUpHorizontalReg_23 ? $signed({{2{_inSpriteX_23_T_4[10]}},_inSpriteX_23_T_4}) :
    $signed(_inSpriteX_23_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1041 = spriteScaleUpHorizontalReg_23 ? _inSpriteHorizontal_23_T_8 : _inSpriteHorizontal_23_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1042 = ~spriteScaleUpHorizontalReg_23 ? $signed({{1{inSpriteXValue_23[11]}},inSpriteXValue_23}) :
    $signed(_GEN_1040); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_23 = ~spriteScaleUpHorizontalReg_23 ? $signed(inSpriteXValue_23) >= 12'sh0 & $signed(
    inSpriteXValue_23) < 12'sh20 : _GEN_1041; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1797 = {{1{spriteYPositionReg_23[9]}},spriteYPositionReg_23}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_23 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1797); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_23 = inSpriteYValue_23[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_23_T = $signed(inSpriteYPreScaled_23) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_23_T_4 = inSpriteYPreScaled_23[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_23_T_8 = _inSpriteVertical_23_T & $signed(inSpriteYPreScaled_23) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_23_T_5 = {$signed(inSpriteYPreScaled_23), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_23_T_14 = _inSpriteVertical_23_T & $signed(inSpriteYPreScaled_23) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1048 = spriteScaleUpVerticalReg_23 ? $signed({{2{_inSpriteY_23_T_4[9]}},_inSpriteY_23_T_4}) :
    $signed(_inSpriteY_23_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1049 = spriteScaleUpVerticalReg_23 ? _inSpriteVertical_23_T_8 : _inSpriteVertical_23_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1050 = ~spriteScaleUpVerticalReg_23 ? $signed({{1{inSpriteYPreScaled_23[10]}},inSpriteYPreScaled_23})
     : $signed(_GEN_1048); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_23 = ~spriteScaleUpVerticalReg_23 ? $signed(inSpriteYPreScaled_23) >= 11'sh0 & $signed(
    inSpriteYPreScaled_23) < 11'sh20 : _GEN_1049; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_24 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_24); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_24_T = $signed(inSpriteXValue_24) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_24_T_4 = inSpriteXValue_24[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_24_T_8 = _inSpriteHorizontal_24_T & $signed(inSpriteXValue_24) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_24_T_5 = {$signed(inSpriteXValue_24), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_24_T_14 = _inSpriteHorizontal_24_T & $signed(inSpriteXValue_24) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1056 = spriteScaleUpHorizontalReg_24 ? $signed({{2{_inSpriteX_24_T_4[10]}},_inSpriteX_24_T_4}) :
    $signed(_inSpriteX_24_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1057 = spriteScaleUpHorizontalReg_24 ? _inSpriteHorizontal_24_T_8 : _inSpriteHorizontal_24_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1058 = ~spriteScaleUpHorizontalReg_24 ? $signed({{1{inSpriteXValue_24[11]}},inSpriteXValue_24}) :
    $signed(_GEN_1056); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_24 = ~spriteScaleUpHorizontalReg_24 ? $signed(inSpriteXValue_24) >= 12'sh0 & $signed(
    inSpriteXValue_24) < 12'sh20 : _GEN_1057; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1799 = {{1{spriteYPositionReg_24[9]}},spriteYPositionReg_24}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_24 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1799); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_24 = inSpriteYValue_24[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_24_T = $signed(inSpriteYPreScaled_24) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_24_T_4 = inSpriteYPreScaled_24[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_24_T_8 = _inSpriteVertical_24_T & $signed(inSpriteYPreScaled_24) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_24_T_5 = {$signed(inSpriteYPreScaled_24), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_24_T_14 = _inSpriteVertical_24_T & $signed(inSpriteYPreScaled_24) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1064 = spriteScaleUpVerticalReg_24 ? $signed({{2{_inSpriteY_24_T_4[9]}},_inSpriteY_24_T_4}) :
    $signed(_inSpriteY_24_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1065 = spriteScaleUpVerticalReg_24 ? _inSpriteVertical_24_T_8 : _inSpriteVertical_24_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1066 = ~spriteScaleUpVerticalReg_24 ? $signed({{1{inSpriteYPreScaled_24[10]}},inSpriteYPreScaled_24})
     : $signed(_GEN_1064); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_24 = ~spriteScaleUpVerticalReg_24 ? $signed(inSpriteYPreScaled_24) >= 11'sh0 & $signed(
    inSpriteYPreScaled_24) < 11'sh20 : _GEN_1065; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_25 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_25); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_25_T = $signed(inSpriteXValue_25) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_25_T_4 = inSpriteXValue_25[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_25_T_8 = _inSpriteHorizontal_25_T & $signed(inSpriteXValue_25) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_25_T_5 = {$signed(inSpriteXValue_25), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_25_T_14 = _inSpriteHorizontal_25_T & $signed(inSpriteXValue_25) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1072 = spriteScaleUpHorizontalReg_25 ? $signed({{2{_inSpriteX_25_T_4[10]}},_inSpriteX_25_T_4}) :
    $signed(_inSpriteX_25_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1073 = spriteScaleUpHorizontalReg_25 ? _inSpriteHorizontal_25_T_8 : _inSpriteHorizontal_25_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1074 = ~spriteScaleUpHorizontalReg_25 ? $signed({{1{inSpriteXValue_25[11]}},inSpriteXValue_25}) :
    $signed(_GEN_1072); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_25 = ~spriteScaleUpHorizontalReg_25 ? $signed(inSpriteXValue_25) >= 12'sh0 & $signed(
    inSpriteXValue_25) < 12'sh20 : _GEN_1073; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1801 = {{1{spriteYPositionReg_25[9]}},spriteYPositionReg_25}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_25 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1801); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_25 = inSpriteYValue_25[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_25_T = $signed(inSpriteYPreScaled_25) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_25_T_4 = inSpriteYPreScaled_25[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_25_T_8 = _inSpriteVertical_25_T & $signed(inSpriteYPreScaled_25) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_25_T_5 = {$signed(inSpriteYPreScaled_25), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_25_T_14 = _inSpriteVertical_25_T & $signed(inSpriteYPreScaled_25) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1080 = spriteScaleUpVerticalReg_25 ? $signed({{2{_inSpriteY_25_T_4[9]}},_inSpriteY_25_T_4}) :
    $signed(_inSpriteY_25_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1081 = spriteScaleUpVerticalReg_25 ? _inSpriteVertical_25_T_8 : _inSpriteVertical_25_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1082 = ~spriteScaleUpVerticalReg_25 ? $signed({{1{inSpriteYPreScaled_25[10]}},inSpriteYPreScaled_25})
     : $signed(_GEN_1080); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_25 = ~spriteScaleUpVerticalReg_25 ? $signed(inSpriteYPreScaled_25) >= 11'sh0 & $signed(
    inSpriteYPreScaled_25) < 11'sh20 : _GEN_1081; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_26 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_26); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_26_T = $signed(inSpriteXValue_26) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_26_T_4 = inSpriteXValue_26[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_26_T_8 = _inSpriteHorizontal_26_T & $signed(inSpriteXValue_26) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_26_T_5 = {$signed(inSpriteXValue_26), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_26_T_14 = _inSpriteHorizontal_26_T & $signed(inSpriteXValue_26) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1088 = spriteScaleUpHorizontalReg_26 ? $signed({{2{_inSpriteX_26_T_4[10]}},_inSpriteX_26_T_4}) :
    $signed(_inSpriteX_26_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1089 = spriteScaleUpHorizontalReg_26 ? _inSpriteHorizontal_26_T_8 : _inSpriteHorizontal_26_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1090 = ~spriteScaleUpHorizontalReg_26 ? $signed({{1{inSpriteXValue_26[11]}},inSpriteXValue_26}) :
    $signed(_GEN_1088); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_26 = ~spriteScaleUpHorizontalReg_26 ? $signed(inSpriteXValue_26) >= 12'sh0 & $signed(
    inSpriteXValue_26) < 12'sh20 : _GEN_1089; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1803 = {{1{spriteYPositionReg_26[9]}},spriteYPositionReg_26}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_26 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1803); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_26 = inSpriteYValue_26[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_26_T = $signed(inSpriteYPreScaled_26) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_26_T_4 = inSpriteYPreScaled_26[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_26_T_8 = _inSpriteVertical_26_T & $signed(inSpriteYPreScaled_26) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_26_T_5 = {$signed(inSpriteYPreScaled_26), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_26_T_14 = _inSpriteVertical_26_T & $signed(inSpriteYPreScaled_26) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1096 = spriteScaleUpVerticalReg_26 ? $signed({{2{_inSpriteY_26_T_4[9]}},_inSpriteY_26_T_4}) :
    $signed(_inSpriteY_26_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1097 = spriteScaleUpVerticalReg_26 ? _inSpriteVertical_26_T_8 : _inSpriteVertical_26_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1098 = ~spriteScaleUpVerticalReg_26 ? $signed({{1{inSpriteYPreScaled_26[10]}},inSpriteYPreScaled_26})
     : $signed(_GEN_1096); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_26 = ~spriteScaleUpVerticalReg_26 ? $signed(inSpriteYPreScaled_26) >= 11'sh0 & $signed(
    inSpriteYPreScaled_26) < 11'sh20 : _GEN_1097; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_27 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_27); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_27_T = $signed(inSpriteXValue_27) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_27_T_4 = inSpriteXValue_27[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_27_T_8 = _inSpriteHorizontal_27_T & $signed(inSpriteXValue_27) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_27_T_5 = {$signed(inSpriteXValue_27), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_27_T_14 = _inSpriteHorizontal_27_T & $signed(inSpriteXValue_27) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1104 = spriteScaleUpHorizontalReg_27 ? $signed({{2{_inSpriteX_27_T_4[10]}},_inSpriteX_27_T_4}) :
    $signed(_inSpriteX_27_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1105 = spriteScaleUpHorizontalReg_27 ? _inSpriteHorizontal_27_T_8 : _inSpriteHorizontal_27_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1106 = ~spriteScaleUpHorizontalReg_27 ? $signed({{1{inSpriteXValue_27[11]}},inSpriteXValue_27}) :
    $signed(_GEN_1104); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_27 = ~spriteScaleUpHorizontalReg_27 ? $signed(inSpriteXValue_27) >= 12'sh0 & $signed(
    inSpriteXValue_27) < 12'sh20 : _GEN_1105; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1805 = {{1{spriteYPositionReg_27[9]}},spriteYPositionReg_27}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_27 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1805); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_27 = inSpriteYValue_27[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_27_T = $signed(inSpriteYPreScaled_27) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_27_T_4 = inSpriteYPreScaled_27[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_27_T_8 = _inSpriteVertical_27_T & $signed(inSpriteYPreScaled_27) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_27_T_5 = {$signed(inSpriteYPreScaled_27), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_27_T_14 = _inSpriteVertical_27_T & $signed(inSpriteYPreScaled_27) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1112 = spriteScaleUpVerticalReg_27 ? $signed({{2{_inSpriteY_27_T_4[9]}},_inSpriteY_27_T_4}) :
    $signed(_inSpriteY_27_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1113 = spriteScaleUpVerticalReg_27 ? _inSpriteVertical_27_T_8 : _inSpriteVertical_27_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1114 = ~spriteScaleUpVerticalReg_27 ? $signed({{1{inSpriteYPreScaled_27[10]}},inSpriteYPreScaled_27})
     : $signed(_GEN_1112); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_27 = ~spriteScaleUpVerticalReg_27 ? $signed(inSpriteYPreScaled_27) >= 11'sh0 & $signed(
    inSpriteYPreScaled_27) < 11'sh20 : _GEN_1113; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_28 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_28); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_28_T = $signed(inSpriteXValue_28) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_28_T_4 = inSpriteXValue_28[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_28_T_8 = _inSpriteHorizontal_28_T & $signed(inSpriteXValue_28) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_28_T_5 = {$signed(inSpriteXValue_28), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_28_T_14 = _inSpriteHorizontal_28_T & $signed(inSpriteXValue_28) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1120 = spriteScaleUpHorizontalReg_28 ? $signed({{2{_inSpriteX_28_T_4[10]}},_inSpriteX_28_T_4}) :
    $signed(_inSpriteX_28_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1121 = spriteScaleUpHorizontalReg_28 ? _inSpriteHorizontal_28_T_8 : _inSpriteHorizontal_28_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1122 = ~spriteScaleUpHorizontalReg_28 ? $signed({{1{inSpriteXValue_28[11]}},inSpriteXValue_28}) :
    $signed(_GEN_1120); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_28 = ~spriteScaleUpHorizontalReg_28 ? $signed(inSpriteXValue_28) >= 12'sh0 & $signed(
    inSpriteXValue_28) < 12'sh20 : _GEN_1121; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1807 = {{1{spriteYPositionReg_28[9]}},spriteYPositionReg_28}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_28 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1807); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_28 = inSpriteYValue_28[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_28_T = $signed(inSpriteYPreScaled_28) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_28_T_4 = inSpriteYPreScaled_28[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_28_T_8 = _inSpriteVertical_28_T & $signed(inSpriteYPreScaled_28) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_28_T_5 = {$signed(inSpriteYPreScaled_28), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_28_T_14 = _inSpriteVertical_28_T & $signed(inSpriteYPreScaled_28) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1128 = spriteScaleUpVerticalReg_28 ? $signed({{2{_inSpriteY_28_T_4[9]}},_inSpriteY_28_T_4}) :
    $signed(_inSpriteY_28_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1129 = spriteScaleUpVerticalReg_28 ? _inSpriteVertical_28_T_8 : _inSpriteVertical_28_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1130 = ~spriteScaleUpVerticalReg_28 ? $signed({{1{inSpriteYPreScaled_28[10]}},inSpriteYPreScaled_28})
     : $signed(_GEN_1128); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_28 = ~spriteScaleUpVerticalReg_28 ? $signed(inSpriteYPreScaled_28) >= 11'sh0 & $signed(
    inSpriteYPreScaled_28) < 11'sh20 : _GEN_1129; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_29 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_29); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_29_T = $signed(inSpriteXValue_29) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_29_T_4 = inSpriteXValue_29[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_29_T_8 = _inSpriteHorizontal_29_T & $signed(inSpriteXValue_29) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_29_T_5 = {$signed(inSpriteXValue_29), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_29_T_14 = _inSpriteHorizontal_29_T & $signed(inSpriteXValue_29) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1136 = spriteScaleUpHorizontalReg_29 ? $signed({{2{_inSpriteX_29_T_4[10]}},_inSpriteX_29_T_4}) :
    $signed(_inSpriteX_29_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1137 = spriteScaleUpHorizontalReg_29 ? _inSpriteHorizontal_29_T_8 : _inSpriteHorizontal_29_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1138 = ~spriteScaleUpHorizontalReg_29 ? $signed({{1{inSpriteXValue_29[11]}},inSpriteXValue_29}) :
    $signed(_GEN_1136); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_29 = ~spriteScaleUpHorizontalReg_29 ? $signed(inSpriteXValue_29) >= 12'sh0 & $signed(
    inSpriteXValue_29) < 12'sh20 : _GEN_1137; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1809 = {{1{spriteYPositionReg_29[9]}},spriteYPositionReg_29}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_29 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1809); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_29 = inSpriteYValue_29[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_29_T = $signed(inSpriteYPreScaled_29) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_29_T_4 = inSpriteYPreScaled_29[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_29_T_8 = _inSpriteVertical_29_T & $signed(inSpriteYPreScaled_29) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_29_T_5 = {$signed(inSpriteYPreScaled_29), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_29_T_14 = _inSpriteVertical_29_T & $signed(inSpriteYPreScaled_29) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1144 = spriteScaleUpVerticalReg_29 ? $signed({{2{_inSpriteY_29_T_4[9]}},_inSpriteY_29_T_4}) :
    $signed(_inSpriteY_29_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1145 = spriteScaleUpVerticalReg_29 ? _inSpriteVertical_29_T_8 : _inSpriteVertical_29_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1146 = ~spriteScaleUpVerticalReg_29 ? $signed({{1{inSpriteYPreScaled_29[10]}},inSpriteYPreScaled_29})
     : $signed(_GEN_1144); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_29 = ~spriteScaleUpVerticalReg_29 ? $signed(inSpriteYPreScaled_29) >= 11'sh0 & $signed(
    inSpriteYPreScaled_29) < 11'sh20 : _GEN_1145; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_30 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_30); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_30_T = $signed(inSpriteXValue_30) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_30_T_4 = inSpriteXValue_30[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_30_T_8 = _inSpriteHorizontal_30_T & $signed(inSpriteXValue_30) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_30_T_5 = {$signed(inSpriteXValue_30), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_30_T_14 = _inSpriteHorizontal_30_T & $signed(inSpriteXValue_30) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1152 = spriteScaleUpHorizontalReg_30 ? $signed({{2{_inSpriteX_30_T_4[10]}},_inSpriteX_30_T_4}) :
    $signed(_inSpriteX_30_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1153 = spriteScaleUpHorizontalReg_30 ? _inSpriteHorizontal_30_T_8 : _inSpriteHorizontal_30_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1154 = ~spriteScaleUpHorizontalReg_30 ? $signed({{1{inSpriteXValue_30[11]}},inSpriteXValue_30}) :
    $signed(_GEN_1152); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_30 = ~spriteScaleUpHorizontalReg_30 ? $signed(inSpriteXValue_30) >= 12'sh0 & $signed(
    inSpriteXValue_30) < 12'sh20 : _GEN_1153; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1811 = {{1{spriteYPositionReg_30[9]}},spriteYPositionReg_30}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_30 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1811); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_30 = inSpriteYValue_30[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_30_T = $signed(inSpriteYPreScaled_30) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_30_T_4 = inSpriteYPreScaled_30[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_30_T_8 = _inSpriteVertical_30_T & $signed(inSpriteYPreScaled_30) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_30_T_5 = {$signed(inSpriteYPreScaled_30), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_30_T_14 = _inSpriteVertical_30_T & $signed(inSpriteYPreScaled_30) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1160 = spriteScaleUpVerticalReg_30 ? $signed({{2{_inSpriteY_30_T_4[9]}},_inSpriteY_30_T_4}) :
    $signed(_inSpriteY_30_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1161 = spriteScaleUpVerticalReg_30 ? _inSpriteVertical_30_T_8 : _inSpriteVertical_30_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1162 = ~spriteScaleUpVerticalReg_30 ? $signed({{1{inSpriteYPreScaled_30[10]}},inSpriteYPreScaled_30})
     : $signed(_GEN_1160); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_30 = ~spriteScaleUpVerticalReg_30 ? $signed(inSpriteYPreScaled_30) >= 11'sh0 & $signed(
    inSpriteYPreScaled_30) < 11'sh20 : _GEN_1161; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_31 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_31); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_31_T = $signed(inSpriteXValue_31) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_31_T_4 = inSpriteXValue_31[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_31_T_8 = _inSpriteHorizontal_31_T & $signed(inSpriteXValue_31) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_31_T_5 = {$signed(inSpriteXValue_31), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_31_T_14 = _inSpriteHorizontal_31_T & $signed(inSpriteXValue_31) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1168 = spriteScaleUpHorizontalReg_31 ? $signed({{2{_inSpriteX_31_T_4[10]}},_inSpriteX_31_T_4}) :
    $signed(_inSpriteX_31_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1169 = spriteScaleUpHorizontalReg_31 ? _inSpriteHorizontal_31_T_8 : _inSpriteHorizontal_31_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1170 = ~spriteScaleUpHorizontalReg_31 ? $signed({{1{inSpriteXValue_31[11]}},inSpriteXValue_31}) :
    $signed(_GEN_1168); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_31 = ~spriteScaleUpHorizontalReg_31 ? $signed(inSpriteXValue_31) >= 12'sh0 & $signed(
    inSpriteXValue_31) < 12'sh20 : _GEN_1169; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1813 = {{1{spriteYPositionReg_31[9]}},spriteYPositionReg_31}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_31 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1813); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_31 = inSpriteYValue_31[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_31_T = $signed(inSpriteYPreScaled_31) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_31_T_4 = inSpriteYPreScaled_31[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_31_T_8 = _inSpriteVertical_31_T & $signed(inSpriteYPreScaled_31) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_31_T_5 = {$signed(inSpriteYPreScaled_31), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_31_T_14 = _inSpriteVertical_31_T & $signed(inSpriteYPreScaled_31) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1176 = spriteScaleUpVerticalReg_31 ? $signed({{2{_inSpriteY_31_T_4[9]}},_inSpriteY_31_T_4}) :
    $signed(_inSpriteY_31_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1177 = spriteScaleUpVerticalReg_31 ? _inSpriteVertical_31_T_8 : _inSpriteVertical_31_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1178 = ~spriteScaleUpVerticalReg_31 ? $signed({{1{inSpriteYPreScaled_31[10]}},inSpriteYPreScaled_31})
     : $signed(_GEN_1176); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_31 = ~spriteScaleUpVerticalReg_31 ? $signed(inSpriteYPreScaled_31) >= 11'sh0 & $signed(
    inSpriteYPreScaled_31) < 11'sh20 : _GEN_1177; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_32 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_32); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_32_T = $signed(inSpriteXValue_32) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_32_T_4 = inSpriteXValue_32[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_32_T_8 = _inSpriteHorizontal_32_T & $signed(inSpriteXValue_32) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_32_T_5 = {$signed(inSpriteXValue_32), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_32_T_14 = _inSpriteHorizontal_32_T & $signed(inSpriteXValue_32) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1184 = spriteScaleUpHorizontalReg_32 ? $signed({{2{_inSpriteX_32_T_4[10]}},_inSpriteX_32_T_4}) :
    $signed(_inSpriteX_32_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1185 = spriteScaleUpHorizontalReg_32 ? _inSpriteHorizontal_32_T_8 : _inSpriteHorizontal_32_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1186 = ~spriteScaleUpHorizontalReg_32 ? $signed({{1{inSpriteXValue_32[11]}},inSpriteXValue_32}) :
    $signed(_GEN_1184); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_32 = ~spriteScaleUpHorizontalReg_32 ? $signed(inSpriteXValue_32) >= 12'sh0 & $signed(
    inSpriteXValue_32) < 12'sh20 : _GEN_1185; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1815 = {{1{spriteYPositionReg_32[9]}},spriteYPositionReg_32}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_32 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1815); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_32 = inSpriteYValue_32[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_32_T = $signed(inSpriteYPreScaled_32) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_32_T_4 = inSpriteYPreScaled_32[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_32_T_8 = _inSpriteVertical_32_T & $signed(inSpriteYPreScaled_32) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_32_T_5 = {$signed(inSpriteYPreScaled_32), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_32_T_14 = _inSpriteVertical_32_T & $signed(inSpriteYPreScaled_32) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1192 = spriteScaleUpVerticalReg_32 ? $signed({{2{_inSpriteY_32_T_4[9]}},_inSpriteY_32_T_4}) :
    $signed(_inSpriteY_32_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1193 = spriteScaleUpVerticalReg_32 ? _inSpriteVertical_32_T_8 : _inSpriteVertical_32_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1194 = ~spriteScaleUpVerticalReg_32 ? $signed({{1{inSpriteYPreScaled_32[10]}},inSpriteYPreScaled_32})
     : $signed(_GEN_1192); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_32 = ~spriteScaleUpVerticalReg_32 ? $signed(inSpriteYPreScaled_32) >= 11'sh0 & $signed(
    inSpriteYPreScaled_32) < 11'sh20 : _GEN_1193; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_33 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_33); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_33_T = $signed(inSpriteXValue_33) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_33_T_4 = inSpriteXValue_33[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_33_T_8 = _inSpriteHorizontal_33_T & $signed(inSpriteXValue_33) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_33_T_5 = {$signed(inSpriteXValue_33), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_33_T_14 = _inSpriteHorizontal_33_T & $signed(inSpriteXValue_33) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1200 = spriteScaleUpHorizontalReg_33 ? $signed({{2{_inSpriteX_33_T_4[10]}},_inSpriteX_33_T_4}) :
    $signed(_inSpriteX_33_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1201 = spriteScaleUpHorizontalReg_33 ? _inSpriteHorizontal_33_T_8 : _inSpriteHorizontal_33_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1202 = ~spriteScaleUpHorizontalReg_33 ? $signed({{1{inSpriteXValue_33[11]}},inSpriteXValue_33}) :
    $signed(_GEN_1200); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_33 = ~spriteScaleUpHorizontalReg_33 ? $signed(inSpriteXValue_33) >= 12'sh0 & $signed(
    inSpriteXValue_33) < 12'sh20 : _GEN_1201; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1817 = {{1{spriteYPositionReg_33[9]}},spriteYPositionReg_33}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_33 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1817); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_33 = inSpriteYValue_33[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_33_T = $signed(inSpriteYPreScaled_33) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_33_T_4 = inSpriteYPreScaled_33[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_33_T_8 = _inSpriteVertical_33_T & $signed(inSpriteYPreScaled_33) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_33_T_5 = {$signed(inSpriteYPreScaled_33), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_33_T_14 = _inSpriteVertical_33_T & $signed(inSpriteYPreScaled_33) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1208 = spriteScaleUpVerticalReg_33 ? $signed({{2{_inSpriteY_33_T_4[9]}},_inSpriteY_33_T_4}) :
    $signed(_inSpriteY_33_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1209 = spriteScaleUpVerticalReg_33 ? _inSpriteVertical_33_T_8 : _inSpriteVertical_33_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1210 = ~spriteScaleUpVerticalReg_33 ? $signed({{1{inSpriteYPreScaled_33[10]}},inSpriteYPreScaled_33})
     : $signed(_GEN_1208); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_33 = ~spriteScaleUpVerticalReg_33 ? $signed(inSpriteYPreScaled_33) >= 11'sh0 & $signed(
    inSpriteYPreScaled_33) < 11'sh20 : _GEN_1209; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_34 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_34); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_34_T = $signed(inSpriteXValue_34) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_34_T_4 = inSpriteXValue_34[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_34_T_8 = _inSpriteHorizontal_34_T & $signed(inSpriteXValue_34) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_34_T_5 = {$signed(inSpriteXValue_34), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_34_T_14 = _inSpriteHorizontal_34_T & $signed(inSpriteXValue_34) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1216 = spriteScaleUpHorizontalReg_34 ? $signed({{2{_inSpriteX_34_T_4[10]}},_inSpriteX_34_T_4}) :
    $signed(_inSpriteX_34_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1217 = spriteScaleUpHorizontalReg_34 ? _inSpriteHorizontal_34_T_8 : _inSpriteHorizontal_34_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1218 = ~spriteScaleUpHorizontalReg_34 ? $signed({{1{inSpriteXValue_34[11]}},inSpriteXValue_34}) :
    $signed(_GEN_1216); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_34 = ~spriteScaleUpHorizontalReg_34 ? $signed(inSpriteXValue_34) >= 12'sh0 & $signed(
    inSpriteXValue_34) < 12'sh20 : _GEN_1217; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1819 = {{1{spriteYPositionReg_34[9]}},spriteYPositionReg_34}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_34 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1819); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_34 = inSpriteYValue_34[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_34_T = $signed(inSpriteYPreScaled_34) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_34_T_4 = inSpriteYPreScaled_34[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_34_T_8 = _inSpriteVertical_34_T & $signed(inSpriteYPreScaled_34) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_34_T_5 = {$signed(inSpriteYPreScaled_34), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_34_T_14 = _inSpriteVertical_34_T & $signed(inSpriteYPreScaled_34) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1224 = spriteScaleUpVerticalReg_34 ? $signed({{2{_inSpriteY_34_T_4[9]}},_inSpriteY_34_T_4}) :
    $signed(_inSpriteY_34_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1225 = spriteScaleUpVerticalReg_34 ? _inSpriteVertical_34_T_8 : _inSpriteVertical_34_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1226 = ~spriteScaleUpVerticalReg_34 ? $signed({{1{inSpriteYPreScaled_34[10]}},inSpriteYPreScaled_34})
     : $signed(_GEN_1224); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_34 = ~spriteScaleUpVerticalReg_34 ? $signed(inSpriteYPreScaled_34) >= 11'sh0 & $signed(
    inSpriteYPreScaled_34) < 11'sh20 : _GEN_1225; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_35 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_35); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_35_T = $signed(inSpriteXValue_35) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_35_T_4 = inSpriteXValue_35[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_35_T_8 = _inSpriteHorizontal_35_T & $signed(inSpriteXValue_35) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_35_T_5 = {$signed(inSpriteXValue_35), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_35_T_14 = _inSpriteHorizontal_35_T & $signed(inSpriteXValue_35) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1232 = spriteScaleUpHorizontalReg_35 ? $signed({{2{_inSpriteX_35_T_4[10]}},_inSpriteX_35_T_4}) :
    $signed(_inSpriteX_35_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1233 = spriteScaleUpHorizontalReg_35 ? _inSpriteHorizontal_35_T_8 : _inSpriteHorizontal_35_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1234 = ~spriteScaleUpHorizontalReg_35 ? $signed({{1{inSpriteXValue_35[11]}},inSpriteXValue_35}) :
    $signed(_GEN_1232); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_35 = ~spriteScaleUpHorizontalReg_35 ? $signed(inSpriteXValue_35) >= 12'sh0 & $signed(
    inSpriteXValue_35) < 12'sh20 : _GEN_1233; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1821 = {{1{spriteYPositionReg_35[9]}},spriteYPositionReg_35}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_35 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1821); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_35 = inSpriteYValue_35[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_35_T = $signed(inSpriteYPreScaled_35) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_35_T_4 = inSpriteYPreScaled_35[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_35_T_8 = _inSpriteVertical_35_T & $signed(inSpriteYPreScaled_35) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_35_T_5 = {$signed(inSpriteYPreScaled_35), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_35_T_14 = _inSpriteVertical_35_T & $signed(inSpriteYPreScaled_35) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1240 = spriteScaleUpVerticalReg_35 ? $signed({{2{_inSpriteY_35_T_4[9]}},_inSpriteY_35_T_4}) :
    $signed(_inSpriteY_35_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1241 = spriteScaleUpVerticalReg_35 ? _inSpriteVertical_35_T_8 : _inSpriteVertical_35_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1242 = ~spriteScaleUpVerticalReg_35 ? $signed({{1{inSpriteYPreScaled_35[10]}},inSpriteYPreScaled_35})
     : $signed(_GEN_1240); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_35 = ~spriteScaleUpVerticalReg_35 ? $signed(inSpriteYPreScaled_35) >= 11'sh0 & $signed(
    inSpriteYPreScaled_35) < 11'sh20 : _GEN_1241; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_36 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_36); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_36_T = $signed(inSpriteXValue_36) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_36_T_4 = inSpriteXValue_36[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_36_T_8 = _inSpriteHorizontal_36_T & $signed(inSpriteXValue_36) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_36_T_5 = {$signed(inSpriteXValue_36), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_36_T_14 = _inSpriteHorizontal_36_T & $signed(inSpriteXValue_36) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1248 = spriteScaleUpHorizontalReg_36 ? $signed({{2{_inSpriteX_36_T_4[10]}},_inSpriteX_36_T_4}) :
    $signed(_inSpriteX_36_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1249 = spriteScaleUpHorizontalReg_36 ? _inSpriteHorizontal_36_T_8 : _inSpriteHorizontal_36_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1250 = ~spriteScaleUpHorizontalReg_36 ? $signed({{1{inSpriteXValue_36[11]}},inSpriteXValue_36}) :
    $signed(_GEN_1248); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_36 = ~spriteScaleUpHorizontalReg_36 ? $signed(inSpriteXValue_36) >= 12'sh0 & $signed(
    inSpriteXValue_36) < 12'sh20 : _GEN_1249; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1823 = {{1{spriteYPositionReg_36[9]}},spriteYPositionReg_36}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_36 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1823); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_36 = inSpriteYValue_36[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_36_T = $signed(inSpriteYPreScaled_36) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_36_T_4 = inSpriteYPreScaled_36[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_36_T_8 = _inSpriteVertical_36_T & $signed(inSpriteYPreScaled_36) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_36_T_5 = {$signed(inSpriteYPreScaled_36), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_36_T_14 = _inSpriteVertical_36_T & $signed(inSpriteYPreScaled_36) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1256 = spriteScaleUpVerticalReg_36 ? $signed({{2{_inSpriteY_36_T_4[9]}},_inSpriteY_36_T_4}) :
    $signed(_inSpriteY_36_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1257 = spriteScaleUpVerticalReg_36 ? _inSpriteVertical_36_T_8 : _inSpriteVertical_36_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1258 = ~spriteScaleUpVerticalReg_36 ? $signed({{1{inSpriteYPreScaled_36[10]}},inSpriteYPreScaled_36})
     : $signed(_GEN_1256); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_36 = ~spriteScaleUpVerticalReg_36 ? $signed(inSpriteYPreScaled_36) >= 11'sh0 & $signed(
    inSpriteYPreScaled_36) < 11'sh20 : _GEN_1257; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_37 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_37); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_37_T = $signed(inSpriteXValue_37) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_37_T_4 = inSpriteXValue_37[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_37_T_8 = _inSpriteHorizontal_37_T & $signed(inSpriteXValue_37) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_37_T_5 = {$signed(inSpriteXValue_37), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_37_T_14 = _inSpriteHorizontal_37_T & $signed(inSpriteXValue_37) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1264 = spriteScaleUpHorizontalReg_37 ? $signed({{2{_inSpriteX_37_T_4[10]}},_inSpriteX_37_T_4}) :
    $signed(_inSpriteX_37_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1265 = spriteScaleUpHorizontalReg_37 ? _inSpriteHorizontal_37_T_8 : _inSpriteHorizontal_37_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1266 = ~spriteScaleUpHorizontalReg_37 ? $signed({{1{inSpriteXValue_37[11]}},inSpriteXValue_37}) :
    $signed(_GEN_1264); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_37 = ~spriteScaleUpHorizontalReg_37 ? $signed(inSpriteXValue_37) >= 12'sh0 & $signed(
    inSpriteXValue_37) < 12'sh20 : _GEN_1265; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1825 = {{1{spriteYPositionReg_37[9]}},spriteYPositionReg_37}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_37 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1825); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_37 = inSpriteYValue_37[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_37_T = $signed(inSpriteYPreScaled_37) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_37_T_4 = inSpriteYPreScaled_37[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_37_T_8 = _inSpriteVertical_37_T & $signed(inSpriteYPreScaled_37) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_37_T_5 = {$signed(inSpriteYPreScaled_37), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_37_T_14 = _inSpriteVertical_37_T & $signed(inSpriteYPreScaled_37) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1272 = spriteScaleUpVerticalReg_37 ? $signed({{2{_inSpriteY_37_T_4[9]}},_inSpriteY_37_T_4}) :
    $signed(_inSpriteY_37_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1273 = spriteScaleUpVerticalReg_37 ? _inSpriteVertical_37_T_8 : _inSpriteVertical_37_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1274 = ~spriteScaleUpVerticalReg_37 ? $signed({{1{inSpriteYPreScaled_37[10]}},inSpriteYPreScaled_37})
     : $signed(_GEN_1272); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_37 = ~spriteScaleUpVerticalReg_37 ? $signed(inSpriteYPreScaled_37) >= 11'sh0 & $signed(
    inSpriteYPreScaled_37) < 11'sh20 : _GEN_1273; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_38 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_38); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_38_T = $signed(inSpriteXValue_38) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_38_T_4 = inSpriteXValue_38[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_38_T_8 = _inSpriteHorizontal_38_T & $signed(inSpriteXValue_38) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_38_T_5 = {$signed(inSpriteXValue_38), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_38_T_14 = _inSpriteHorizontal_38_T & $signed(inSpriteXValue_38) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1280 = spriteScaleUpHorizontalReg_38 ? $signed({{2{_inSpriteX_38_T_4[10]}},_inSpriteX_38_T_4}) :
    $signed(_inSpriteX_38_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1281 = spriteScaleUpHorizontalReg_38 ? _inSpriteHorizontal_38_T_8 : _inSpriteHorizontal_38_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1282 = ~spriteScaleUpHorizontalReg_38 ? $signed({{1{inSpriteXValue_38[11]}},inSpriteXValue_38}) :
    $signed(_GEN_1280); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_38 = ~spriteScaleUpHorizontalReg_38 ? $signed(inSpriteXValue_38) >= 12'sh0 & $signed(
    inSpriteXValue_38) < 12'sh20 : _GEN_1281; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1827 = {{1{spriteYPositionReg_38[9]}},spriteYPositionReg_38}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_38 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1827); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_38 = inSpriteYValue_38[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_38_T = $signed(inSpriteYPreScaled_38) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_38_T_4 = inSpriteYPreScaled_38[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_38_T_8 = _inSpriteVertical_38_T & $signed(inSpriteYPreScaled_38) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_38_T_5 = {$signed(inSpriteYPreScaled_38), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_38_T_14 = _inSpriteVertical_38_T & $signed(inSpriteYPreScaled_38) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1288 = spriteScaleUpVerticalReg_38 ? $signed({{2{_inSpriteY_38_T_4[9]}},_inSpriteY_38_T_4}) :
    $signed(_inSpriteY_38_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1289 = spriteScaleUpVerticalReg_38 ? _inSpriteVertical_38_T_8 : _inSpriteVertical_38_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1290 = ~spriteScaleUpVerticalReg_38 ? $signed({{1{inSpriteYPreScaled_38[10]}},inSpriteYPreScaled_38})
     : $signed(_GEN_1288); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_38 = ~spriteScaleUpVerticalReg_38 ? $signed(inSpriteYPreScaled_38) >= 11'sh0 & $signed(
    inSpriteYPreScaled_38) < 11'sh20 : _GEN_1289; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_39 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_39); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_39_T = $signed(inSpriteXValue_39) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_39_T_4 = inSpriteXValue_39[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_39_T_8 = _inSpriteHorizontal_39_T & $signed(inSpriteXValue_39) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_39_T_5 = {$signed(inSpriteXValue_39), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_39_T_14 = _inSpriteHorizontal_39_T & $signed(inSpriteXValue_39) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1296 = spriteScaleUpHorizontalReg_39 ? $signed({{2{_inSpriteX_39_T_4[10]}},_inSpriteX_39_T_4}) :
    $signed(_inSpriteX_39_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1297 = spriteScaleUpHorizontalReg_39 ? _inSpriteHorizontal_39_T_8 : _inSpriteHorizontal_39_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1298 = ~spriteScaleUpHorizontalReg_39 ? $signed({{1{inSpriteXValue_39[11]}},inSpriteXValue_39}) :
    $signed(_GEN_1296); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_39 = ~spriteScaleUpHorizontalReg_39 ? $signed(inSpriteXValue_39) >= 12'sh0 & $signed(
    inSpriteXValue_39) < 12'sh20 : _GEN_1297; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1829 = {{1{spriteYPositionReg_39[9]}},spriteYPositionReg_39}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_39 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1829); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_39 = inSpriteYValue_39[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_39_T = $signed(inSpriteYPreScaled_39) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_39_T_4 = inSpriteYPreScaled_39[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_39_T_8 = _inSpriteVertical_39_T & $signed(inSpriteYPreScaled_39) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_39_T_5 = {$signed(inSpriteYPreScaled_39), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_39_T_14 = _inSpriteVertical_39_T & $signed(inSpriteYPreScaled_39) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1304 = spriteScaleUpVerticalReg_39 ? $signed({{2{_inSpriteY_39_T_4[9]}},_inSpriteY_39_T_4}) :
    $signed(_inSpriteY_39_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1305 = spriteScaleUpVerticalReg_39 ? _inSpriteVertical_39_T_8 : _inSpriteVertical_39_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1306 = ~spriteScaleUpVerticalReg_39 ? $signed({{1{inSpriteYPreScaled_39[10]}},inSpriteYPreScaled_39})
     : $signed(_GEN_1304); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_39 = ~spriteScaleUpVerticalReg_39 ? $signed(inSpriteYPreScaled_39) >= 11'sh0 & $signed(
    inSpriteYPreScaled_39) < 11'sh20 : _GEN_1305; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_40 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_40); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_40_T = $signed(inSpriteXValue_40) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_40_T_4 = inSpriteXValue_40[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_40_T_8 = _inSpriteHorizontal_40_T & $signed(inSpriteXValue_40) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_40_T_5 = {$signed(inSpriteXValue_40), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_40_T_14 = _inSpriteHorizontal_40_T & $signed(inSpriteXValue_40) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1312 = spriteScaleUpHorizontalReg_40 ? $signed({{2{_inSpriteX_40_T_4[10]}},_inSpriteX_40_T_4}) :
    $signed(_inSpriteX_40_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1313 = spriteScaleUpHorizontalReg_40 ? _inSpriteHorizontal_40_T_8 : _inSpriteHorizontal_40_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1314 = ~spriteScaleUpHorizontalReg_40 ? $signed({{1{inSpriteXValue_40[11]}},inSpriteXValue_40}) :
    $signed(_GEN_1312); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_40 = ~spriteScaleUpHorizontalReg_40 ? $signed(inSpriteXValue_40) >= 12'sh0 & $signed(
    inSpriteXValue_40) < 12'sh20 : _GEN_1313; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1831 = {{1{spriteYPositionReg_40[9]}},spriteYPositionReg_40}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_40 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1831); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_40 = inSpriteYValue_40[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_40_T = $signed(inSpriteYPreScaled_40) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_40_T_4 = inSpriteYPreScaled_40[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_40_T_8 = _inSpriteVertical_40_T & $signed(inSpriteYPreScaled_40) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_40_T_5 = {$signed(inSpriteYPreScaled_40), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_40_T_14 = _inSpriteVertical_40_T & $signed(inSpriteYPreScaled_40) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1320 = spriteScaleUpVerticalReg_40 ? $signed({{2{_inSpriteY_40_T_4[9]}},_inSpriteY_40_T_4}) :
    $signed(_inSpriteY_40_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1321 = spriteScaleUpVerticalReg_40 ? _inSpriteVertical_40_T_8 : _inSpriteVertical_40_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1322 = ~spriteScaleUpVerticalReg_40 ? $signed({{1{inSpriteYPreScaled_40[10]}},inSpriteYPreScaled_40})
     : $signed(_GEN_1320); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_40 = ~spriteScaleUpVerticalReg_40 ? $signed(inSpriteYPreScaled_40) >= 11'sh0 & $signed(
    inSpriteYPreScaled_40) < 11'sh20 : _GEN_1321; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_41 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_41); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_41_T = $signed(inSpriteXValue_41) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_41_T_4 = inSpriteXValue_41[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_41_T_8 = _inSpriteHorizontal_41_T & $signed(inSpriteXValue_41) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_41_T_5 = {$signed(inSpriteXValue_41), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_41_T_14 = _inSpriteHorizontal_41_T & $signed(inSpriteXValue_41) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1328 = spriteScaleUpHorizontalReg_41 ? $signed({{2{_inSpriteX_41_T_4[10]}},_inSpriteX_41_T_4}) :
    $signed(_inSpriteX_41_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1329 = spriteScaleUpHorizontalReg_41 ? _inSpriteHorizontal_41_T_8 : _inSpriteHorizontal_41_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1330 = ~spriteScaleUpHorizontalReg_41 ? $signed({{1{inSpriteXValue_41[11]}},inSpriteXValue_41}) :
    $signed(_GEN_1328); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_41 = ~spriteScaleUpHorizontalReg_41 ? $signed(inSpriteXValue_41) >= 12'sh0 & $signed(
    inSpriteXValue_41) < 12'sh20 : _GEN_1329; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1833 = {{1{spriteYPositionReg_41[9]}},spriteYPositionReg_41}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_41 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1833); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_41 = inSpriteYValue_41[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_41_T = $signed(inSpriteYPreScaled_41) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_41_T_4 = inSpriteYPreScaled_41[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_41_T_8 = _inSpriteVertical_41_T & $signed(inSpriteYPreScaled_41) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_41_T_5 = {$signed(inSpriteYPreScaled_41), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_41_T_14 = _inSpriteVertical_41_T & $signed(inSpriteYPreScaled_41) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1336 = spriteScaleUpVerticalReg_41 ? $signed({{2{_inSpriteY_41_T_4[9]}},_inSpriteY_41_T_4}) :
    $signed(_inSpriteY_41_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1337 = spriteScaleUpVerticalReg_41 ? _inSpriteVertical_41_T_8 : _inSpriteVertical_41_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1338 = ~spriteScaleUpVerticalReg_41 ? $signed({{1{inSpriteYPreScaled_41[10]}},inSpriteYPreScaled_41})
     : $signed(_GEN_1336); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_41 = ~spriteScaleUpVerticalReg_41 ? $signed(inSpriteYPreScaled_41) >= 11'sh0 & $signed(
    inSpriteYPreScaled_41) < 11'sh20 : _GEN_1337; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_42 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_42); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_42_T = $signed(inSpriteXValue_42) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_42_T_4 = inSpriteXValue_42[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_42_T_8 = _inSpriteHorizontal_42_T & $signed(inSpriteXValue_42) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_42_T_5 = {$signed(inSpriteXValue_42), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_42_T_14 = _inSpriteHorizontal_42_T & $signed(inSpriteXValue_42) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1344 = spriteScaleUpHorizontalReg_42 ? $signed({{2{_inSpriteX_42_T_4[10]}},_inSpriteX_42_T_4}) :
    $signed(_inSpriteX_42_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1345 = spriteScaleUpHorizontalReg_42 ? _inSpriteHorizontal_42_T_8 : _inSpriteHorizontal_42_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1346 = ~spriteScaleUpHorizontalReg_42 ? $signed({{1{inSpriteXValue_42[11]}},inSpriteXValue_42}) :
    $signed(_GEN_1344); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_42 = ~spriteScaleUpHorizontalReg_42 ? $signed(inSpriteXValue_42) >= 12'sh0 & $signed(
    inSpriteXValue_42) < 12'sh20 : _GEN_1345; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1835 = {{1{spriteYPositionReg_42[9]}},spriteYPositionReg_42}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_42 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1835); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_42 = inSpriteYValue_42[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_42_T = $signed(inSpriteYPreScaled_42) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_42_T_4 = inSpriteYPreScaled_42[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_42_T_8 = _inSpriteVertical_42_T & $signed(inSpriteYPreScaled_42) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_42_T_5 = {$signed(inSpriteYPreScaled_42), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_42_T_14 = _inSpriteVertical_42_T & $signed(inSpriteYPreScaled_42) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1352 = spriteScaleUpVerticalReg_42 ? $signed({{2{_inSpriteY_42_T_4[9]}},_inSpriteY_42_T_4}) :
    $signed(_inSpriteY_42_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1353 = spriteScaleUpVerticalReg_42 ? _inSpriteVertical_42_T_8 : _inSpriteVertical_42_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1354 = ~spriteScaleUpVerticalReg_42 ? $signed({{1{inSpriteYPreScaled_42[10]}},inSpriteYPreScaled_42})
     : $signed(_GEN_1352); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_42 = ~spriteScaleUpVerticalReg_42 ? $signed(inSpriteYPreScaled_42) >= 11'sh0 & $signed(
    inSpriteYPreScaled_42) < 11'sh20 : _GEN_1353; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_43 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_43); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_43_T = $signed(inSpriteXValue_43) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_43_T_4 = inSpriteXValue_43[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_43_T_8 = _inSpriteHorizontal_43_T & $signed(inSpriteXValue_43) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_43_T_5 = {$signed(inSpriteXValue_43), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_43_T_14 = _inSpriteHorizontal_43_T & $signed(inSpriteXValue_43) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1360 = spriteScaleUpHorizontalReg_43 ? $signed({{2{_inSpriteX_43_T_4[10]}},_inSpriteX_43_T_4}) :
    $signed(_inSpriteX_43_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1361 = spriteScaleUpHorizontalReg_43 ? _inSpriteHorizontal_43_T_8 : _inSpriteHorizontal_43_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1362 = ~spriteScaleUpHorizontalReg_43 ? $signed({{1{inSpriteXValue_43[11]}},inSpriteXValue_43}) :
    $signed(_GEN_1360); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_43 = ~spriteScaleUpHorizontalReg_43 ? $signed(inSpriteXValue_43) >= 12'sh0 & $signed(
    inSpriteXValue_43) < 12'sh20 : _GEN_1361; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1837 = {{1{spriteYPositionReg_43[9]}},spriteYPositionReg_43}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_43 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1837); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_43 = inSpriteYValue_43[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_43_T = $signed(inSpriteYPreScaled_43) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_43_T_4 = inSpriteYPreScaled_43[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_43_T_8 = _inSpriteVertical_43_T & $signed(inSpriteYPreScaled_43) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_43_T_5 = {$signed(inSpriteYPreScaled_43), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_43_T_14 = _inSpriteVertical_43_T & $signed(inSpriteYPreScaled_43) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1368 = spriteScaleUpVerticalReg_43 ? $signed({{2{_inSpriteY_43_T_4[9]}},_inSpriteY_43_T_4}) :
    $signed(_inSpriteY_43_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1369 = spriteScaleUpVerticalReg_43 ? _inSpriteVertical_43_T_8 : _inSpriteVertical_43_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1370 = ~spriteScaleUpVerticalReg_43 ? $signed({{1{inSpriteYPreScaled_43[10]}},inSpriteYPreScaled_43})
     : $signed(_GEN_1368); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_43 = ~spriteScaleUpVerticalReg_43 ? $signed(inSpriteYPreScaled_43) >= 11'sh0 & $signed(
    inSpriteYPreScaled_43) < 11'sh20 : _GEN_1369; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_44 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_44); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_44_T = $signed(inSpriteXValue_44) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_44_T_4 = inSpriteXValue_44[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_44_T_8 = _inSpriteHorizontal_44_T & $signed(inSpriteXValue_44) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_44_T_5 = {$signed(inSpriteXValue_44), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_44_T_14 = _inSpriteHorizontal_44_T & $signed(inSpriteXValue_44) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1376 = spriteScaleUpHorizontalReg_44 ? $signed({{2{_inSpriteX_44_T_4[10]}},_inSpriteX_44_T_4}) :
    $signed(_inSpriteX_44_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1377 = spriteScaleUpHorizontalReg_44 ? _inSpriteHorizontal_44_T_8 : _inSpriteHorizontal_44_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1378 = ~spriteScaleUpHorizontalReg_44 ? $signed({{1{inSpriteXValue_44[11]}},inSpriteXValue_44}) :
    $signed(_GEN_1376); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_44 = ~spriteScaleUpHorizontalReg_44 ? $signed(inSpriteXValue_44) >= 12'sh0 & $signed(
    inSpriteXValue_44) < 12'sh20 : _GEN_1377; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1839 = {{1{spriteYPositionReg_44[9]}},spriteYPositionReg_44}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_44 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1839); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_44 = inSpriteYValue_44[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_44_T = $signed(inSpriteYPreScaled_44) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_44_T_4 = inSpriteYPreScaled_44[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_44_T_8 = _inSpriteVertical_44_T & $signed(inSpriteYPreScaled_44) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_44_T_5 = {$signed(inSpriteYPreScaled_44), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_44_T_14 = _inSpriteVertical_44_T & $signed(inSpriteYPreScaled_44) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1384 = spriteScaleUpVerticalReg_44 ? $signed({{2{_inSpriteY_44_T_4[9]}},_inSpriteY_44_T_4}) :
    $signed(_inSpriteY_44_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1385 = spriteScaleUpVerticalReg_44 ? _inSpriteVertical_44_T_8 : _inSpriteVertical_44_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1386 = ~spriteScaleUpVerticalReg_44 ? $signed({{1{inSpriteYPreScaled_44[10]}},inSpriteYPreScaled_44})
     : $signed(_GEN_1384); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_44 = ~spriteScaleUpVerticalReg_44 ? $signed(inSpriteYPreScaled_44) >= 11'sh0 & $signed(
    inSpriteYPreScaled_44) < 11'sh20 : _GEN_1385; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_45 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_45); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_45_T = $signed(inSpriteXValue_45) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_45_T_4 = inSpriteXValue_45[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_45_T_8 = _inSpriteHorizontal_45_T & $signed(inSpriteXValue_45) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_45_T_5 = {$signed(inSpriteXValue_45), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_45_T_14 = _inSpriteHorizontal_45_T & $signed(inSpriteXValue_45) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1392 = spriteScaleUpHorizontalReg_45 ? $signed({{2{_inSpriteX_45_T_4[10]}},_inSpriteX_45_T_4}) :
    $signed(_inSpriteX_45_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1393 = spriteScaleUpHorizontalReg_45 ? _inSpriteHorizontal_45_T_8 : _inSpriteHorizontal_45_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1394 = ~spriteScaleUpHorizontalReg_45 ? $signed({{1{inSpriteXValue_45[11]}},inSpriteXValue_45}) :
    $signed(_GEN_1392); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_45 = ~spriteScaleUpHorizontalReg_45 ? $signed(inSpriteXValue_45) >= 12'sh0 & $signed(
    inSpriteXValue_45) < 12'sh20 : _GEN_1393; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1841 = {{1{spriteYPositionReg_45[9]}},spriteYPositionReg_45}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_45 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1841); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_45 = inSpriteYValue_45[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_45_T = $signed(inSpriteYPreScaled_45) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_45_T_4 = inSpriteYPreScaled_45[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_45_T_8 = _inSpriteVertical_45_T & $signed(inSpriteYPreScaled_45) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_45_T_5 = {$signed(inSpriteYPreScaled_45), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_45_T_14 = _inSpriteVertical_45_T & $signed(inSpriteYPreScaled_45) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1400 = spriteScaleUpVerticalReg_45 ? $signed({{2{_inSpriteY_45_T_4[9]}},_inSpriteY_45_T_4}) :
    $signed(_inSpriteY_45_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1401 = spriteScaleUpVerticalReg_45 ? _inSpriteVertical_45_T_8 : _inSpriteVertical_45_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1402 = ~spriteScaleUpVerticalReg_45 ? $signed({{1{inSpriteYPreScaled_45[10]}},inSpriteYPreScaled_45})
     : $signed(_GEN_1400); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_45 = ~spriteScaleUpVerticalReg_45 ? $signed(inSpriteYPreScaled_45) >= 11'sh0 & $signed(
    inSpriteYPreScaled_45) < 11'sh20 : _GEN_1401; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_46 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_46); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_46 = $signed(inSpriteXValue_46) >= 12'sh0 & $signed(inSpriteXValue_46) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1410 = {{1{inSpriteXValue_46[11]}},inSpriteXValue_46}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1843 = {{1{spriteYPositionReg_46[9]}},spriteYPositionReg_46}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_46 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1843); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_46 = inSpriteYValue_46[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_46 = $signed(inSpriteYPreScaled_46) >= 11'sh0 & $signed(inSpriteYPreScaled_46) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1418 = {{1{inSpriteYPreScaled_46[10]}},inSpriteYPreScaled_46}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_47 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_47); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_47 = $signed(inSpriteXValue_47) >= 12'sh0 & $signed(inSpriteXValue_47) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1426 = {{1{inSpriteXValue_47[11]}},inSpriteXValue_47}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1845 = {{1{spriteYPositionReg_47[9]}},spriteYPositionReg_47}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_47 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1845); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_47 = inSpriteYValue_47[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_47 = $signed(inSpriteYPreScaled_47) >= 11'sh0 & $signed(inSpriteYPreScaled_47) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1434 = {{1{inSpriteYPreScaled_47[10]}},inSpriteYPreScaled_47}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_48 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_48); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_48 = $signed(inSpriteXValue_48) >= 12'sh0 & $signed(inSpriteXValue_48) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1442 = {{1{inSpriteXValue_48[11]}},inSpriteXValue_48}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1847 = {{1{spriteYPositionReg_48[9]}},spriteYPositionReg_48}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_48 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1847); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_48 = inSpriteYValue_48[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_48 = $signed(inSpriteYPreScaled_48) >= 11'sh0 & $signed(inSpriteYPreScaled_48) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1450 = {{1{inSpriteYPreScaled_48[10]}},inSpriteYPreScaled_48}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_49 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_49); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_49 = $signed(inSpriteXValue_49) >= 12'sh0 & $signed(inSpriteXValue_49) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1458 = {{1{inSpriteXValue_49[11]}},inSpriteXValue_49}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1849 = {{1{spriteYPositionReg_49[9]}},spriteYPositionReg_49}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_49 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1849); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_49 = inSpriteYValue_49[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_49 = $signed(inSpriteYPreScaled_49) >= 11'sh0 & $signed(inSpriteYPreScaled_49) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1466 = {{1{inSpriteYPreScaled_49[10]}},inSpriteYPreScaled_49}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_50 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_50); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_50 = $signed(inSpriteXValue_50) >= 12'sh0 & $signed(inSpriteXValue_50) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1474 = {{1{inSpriteXValue_50[11]}},inSpriteXValue_50}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1851 = {{1{spriteYPositionReg_50[9]}},spriteYPositionReg_50}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_50 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1851); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_50 = inSpriteYValue_50[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_50 = $signed(inSpriteYPreScaled_50) >= 11'sh0 & $signed(inSpriteYPreScaled_50) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1482 = {{1{inSpriteYPreScaled_50[10]}},inSpriteYPreScaled_50}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_51 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_51); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_51 = $signed(inSpriteXValue_51) >= 12'sh0 & $signed(inSpriteXValue_51) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1490 = {{1{inSpriteXValue_51[11]}},inSpriteXValue_51}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1853 = {{1{spriteYPositionReg_51[9]}},spriteYPositionReg_51}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_51 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1853); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_51 = inSpriteYValue_51[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_51 = $signed(inSpriteYPreScaled_51) >= 11'sh0 & $signed(inSpriteYPreScaled_51) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1498 = {{1{inSpriteYPreScaled_51[10]}},inSpriteYPreScaled_51}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_52 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_52); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_52 = $signed(inSpriteXValue_52) >= 12'sh0 & $signed(inSpriteXValue_52) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1506 = {{1{inSpriteXValue_52[11]}},inSpriteXValue_52}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1855 = {{1{spriteYPositionReg_52[9]}},spriteYPositionReg_52}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_52 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1855); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_52 = inSpriteYValue_52[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_52 = $signed(inSpriteYPreScaled_52) >= 11'sh0 & $signed(inSpriteYPreScaled_52) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1514 = {{1{inSpriteYPreScaled_52[10]}},inSpriteYPreScaled_52}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_53 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_53); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_53 = $signed(inSpriteXValue_53) >= 12'sh0 & $signed(inSpriteXValue_53) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1522 = {{1{inSpriteXValue_53[11]}},inSpriteXValue_53}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1857 = {{1{spriteYPositionReg_53[9]}},spriteYPositionReg_53}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_53 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1857); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_53 = inSpriteYValue_53[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_53 = $signed(inSpriteYPreScaled_53) >= 11'sh0 & $signed(inSpriteYPreScaled_53) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1530 = {{1{inSpriteYPreScaled_53[10]}},inSpriteYPreScaled_53}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_54 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_54); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_54 = $signed(inSpriteXValue_54) >= 12'sh0 & $signed(inSpriteXValue_54) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1538 = {{1{inSpriteXValue_54[11]}},inSpriteXValue_54}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1859 = {{1{spriteYPositionReg_54[9]}},spriteYPositionReg_54}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_54 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1859); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_54 = inSpriteYValue_54[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_54 = $signed(inSpriteYPreScaled_54) >= 11'sh0 & $signed(inSpriteYPreScaled_54) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1546 = {{1{inSpriteYPreScaled_54[10]}},inSpriteYPreScaled_54}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_55 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_55); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_55 = $signed(inSpriteXValue_55) >= 12'sh0 & $signed(inSpriteXValue_55) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1554 = {{1{inSpriteXValue_55[11]}},inSpriteXValue_55}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1861 = {{1{spriteYPositionReg_55[9]}},spriteYPositionReg_55}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_55 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1861); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_55 = inSpriteYValue_55[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_55 = $signed(inSpriteYPreScaled_55) >= 11'sh0 & $signed(inSpriteYPreScaled_55) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1562 = {{1{inSpriteYPreScaled_55[10]}},inSpriteYPreScaled_55}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_56 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_56); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_56 = $signed(inSpriteXValue_56) >= 12'sh0 & $signed(inSpriteXValue_56) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1570 = {{1{inSpriteXValue_56[11]}},inSpriteXValue_56}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1863 = {{1{spriteYPositionReg_56[9]}},spriteYPositionReg_56}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_56 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1863); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_56 = inSpriteYValue_56[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_56 = $signed(inSpriteYPreScaled_56) >= 11'sh0 & $signed(inSpriteYPreScaled_56) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1578 = {{1{inSpriteYPreScaled_56[10]}},inSpriteYPreScaled_56}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_57 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_57); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_57 = $signed(inSpriteXValue_57) >= 12'sh0 & $signed(inSpriteXValue_57) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1586 = {{1{inSpriteXValue_57[11]}},inSpriteXValue_57}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1865 = {{1{spriteYPositionReg_57[9]}},spriteYPositionReg_57}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_57 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1865); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_57 = inSpriteYValue_57[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_57 = $signed(inSpriteYPreScaled_57) >= 11'sh0 & $signed(inSpriteYPreScaled_57) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1594 = {{1{inSpriteYPreScaled_57[10]}},inSpriteYPreScaled_57}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_58 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_58); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_58_T = $signed(inSpriteXValue_58) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_58_T_4 = inSpriteXValue_58[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_58_T_8 = _inSpriteHorizontal_58_T & $signed(inSpriteXValue_58) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_58_T_5 = {$signed(inSpriteXValue_58), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_58_T_14 = _inSpriteHorizontal_58_T & $signed(inSpriteXValue_58) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1600 = spriteScaleUpHorizontalReg_58 ? $signed({{2{_inSpriteX_58_T_4[10]}},_inSpriteX_58_T_4}) :
    $signed(_inSpriteX_58_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1601 = spriteScaleUpHorizontalReg_58 ? _inSpriteHorizontal_58_T_8 : _inSpriteHorizontal_58_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1602 = ~spriteScaleUpHorizontalReg_58 ? $signed({{1{inSpriteXValue_58[11]}},inSpriteXValue_58}) :
    $signed(_GEN_1600); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_58 = ~spriteScaleUpHorizontalReg_58 ? $signed(inSpriteXValue_58) >= 12'sh0 & $signed(
    inSpriteXValue_58) < 12'sh20 : _GEN_1601; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1867 = {{1{spriteYPositionReg_58[9]}},spriteYPositionReg_58}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_58 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1867); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_58 = inSpriteYValue_58[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_58_T = $signed(inSpriteYPreScaled_58) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_58_T_4 = inSpriteYPreScaled_58[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_58_T_8 = _inSpriteVertical_58_T & $signed(inSpriteYPreScaled_58) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_58_T_5 = {$signed(inSpriteYPreScaled_58), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_58_T_14 = _inSpriteVertical_58_T & $signed(inSpriteYPreScaled_58) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1608 = spriteScaleUpVerticalReg_58 ? $signed({{2{_inSpriteY_58_T_4[9]}},_inSpriteY_58_T_4}) :
    $signed(_inSpriteY_58_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1609 = spriteScaleUpVerticalReg_58 ? _inSpriteVertical_58_T_8 : _inSpriteVertical_58_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1610 = ~spriteScaleUpVerticalReg_58 ? $signed({{1{inSpriteYPreScaled_58[10]}},inSpriteYPreScaled_58})
     : $signed(_GEN_1608); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_58 = ~spriteScaleUpVerticalReg_58 ? $signed(inSpriteYPreScaled_58) >= 11'sh0 & $signed(
    inSpriteYPreScaled_58) < 11'sh20 : _GEN_1609; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_59 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_59); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_59_T = $signed(inSpriteXValue_59) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_59_T_4 = inSpriteXValue_59[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_59_T_8 = _inSpriteHorizontal_59_T & $signed(inSpriteXValue_59) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_59_T_5 = {$signed(inSpriteXValue_59), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_59_T_14 = _inSpriteHorizontal_59_T & $signed(inSpriteXValue_59) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1616 = spriteScaleUpHorizontalReg_59 ? $signed({{2{_inSpriteX_59_T_4[10]}},_inSpriteX_59_T_4}) :
    $signed(_inSpriteX_59_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1617 = spriteScaleUpHorizontalReg_59 ? _inSpriteHorizontal_59_T_8 : _inSpriteHorizontal_59_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1618 = ~spriteScaleUpHorizontalReg_59 ? $signed({{1{inSpriteXValue_59[11]}},inSpriteXValue_59}) :
    $signed(_GEN_1616); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_59 = ~spriteScaleUpHorizontalReg_59 ? $signed(inSpriteXValue_59) >= 12'sh0 & $signed(
    inSpriteXValue_59) < 12'sh20 : _GEN_1617; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1869 = {{1{spriteYPositionReg_59[9]}},spriteYPositionReg_59}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_59 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1869); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_59 = inSpriteYValue_59[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_59_T = $signed(inSpriteYPreScaled_59) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_59_T_4 = inSpriteYPreScaled_59[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_59_T_8 = _inSpriteVertical_59_T & $signed(inSpriteYPreScaled_59) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_59_T_5 = {$signed(inSpriteYPreScaled_59), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_59_T_14 = _inSpriteVertical_59_T & $signed(inSpriteYPreScaled_59) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1624 = spriteScaleUpVerticalReg_59 ? $signed({{2{_inSpriteY_59_T_4[9]}},_inSpriteY_59_T_4}) :
    $signed(_inSpriteY_59_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1625 = spriteScaleUpVerticalReg_59 ? _inSpriteVertical_59_T_8 : _inSpriteVertical_59_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1626 = ~spriteScaleUpVerticalReg_59 ? $signed({{1{inSpriteYPreScaled_59[10]}},inSpriteYPreScaled_59})
     : $signed(_GEN_1624); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_59 = ~spriteScaleUpVerticalReg_59 ? $signed(inSpriteYPreScaled_59) >= 11'sh0 & $signed(
    inSpriteYPreScaled_59) < 11'sh20 : _GEN_1625; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_60 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_60); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_60_T = $signed(inSpriteXValue_60) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_60_T_4 = inSpriteXValue_60[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_60_T_8 = _inSpriteHorizontal_60_T & $signed(inSpriteXValue_60) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_60_T_5 = {$signed(inSpriteXValue_60), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_60_T_14 = _inSpriteHorizontal_60_T & $signed(inSpriteXValue_60) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1632 = spriteScaleUpHorizontalReg_60 ? $signed({{2{_inSpriteX_60_T_4[10]}},_inSpriteX_60_T_4}) :
    $signed(_inSpriteX_60_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1633 = spriteScaleUpHorizontalReg_60 ? _inSpriteHorizontal_60_T_8 : _inSpriteHorizontal_60_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1634 = ~spriteScaleUpHorizontalReg_60 ? $signed({{1{inSpriteXValue_60[11]}},inSpriteXValue_60}) :
    $signed(_GEN_1632); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_60 = ~spriteScaleUpHorizontalReg_60 ? $signed(inSpriteXValue_60) >= 12'sh0 & $signed(
    inSpriteXValue_60) < 12'sh20 : _GEN_1633; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1871 = {{1{spriteYPositionReg_60[9]}},spriteYPositionReg_60}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_60 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1871); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_60 = inSpriteYValue_60[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_60_T = $signed(inSpriteYPreScaled_60) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_60_T_4 = inSpriteYPreScaled_60[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_60_T_8 = _inSpriteVertical_60_T & $signed(inSpriteYPreScaled_60) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_60_T_5 = {$signed(inSpriteYPreScaled_60), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_60_T_14 = _inSpriteVertical_60_T & $signed(inSpriteYPreScaled_60) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1640 = spriteScaleUpVerticalReg_60 ? $signed({{2{_inSpriteY_60_T_4[9]}},_inSpriteY_60_T_4}) :
    $signed(_inSpriteY_60_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1641 = spriteScaleUpVerticalReg_60 ? _inSpriteVertical_60_T_8 : _inSpriteVertical_60_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1642 = ~spriteScaleUpVerticalReg_60 ? $signed({{1{inSpriteYPreScaled_60[10]}},inSpriteYPreScaled_60})
     : $signed(_GEN_1640); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_60 = ~spriteScaleUpVerticalReg_60 ? $signed(inSpriteYPreScaled_60) >= 11'sh0 & $signed(
    inSpriteYPreScaled_60) < 11'sh20 : _GEN_1641; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_61 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_61); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_61 = $signed(inSpriteXValue_61) >= 12'sh0 & $signed(inSpriteXValue_61) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1650 = {{1{inSpriteXValue_61[11]}},inSpriteXValue_61}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1873 = {{1{spriteYPositionReg_61[9]}},spriteYPositionReg_61}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_61 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1873); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_61 = inSpriteYValue_61[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_61 = $signed(inSpriteYPreScaled_61) >= 11'sh0 & $signed(inSpriteYPreScaled_61) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1658 = {{1{inSpriteYPreScaled_61[10]}},inSpriteYPreScaled_61}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_62 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_62); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_62 = $signed(inSpriteXValue_62) >= 12'sh0 & $signed(inSpriteXValue_62) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1666 = {{1{inSpriteXValue_62[11]}},inSpriteXValue_62}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1875 = {{1{spriteYPositionReg_62[9]}},spriteYPositionReg_62}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_62 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1875); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_62 = inSpriteYValue_62[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_62 = $signed(inSpriteYPreScaled_62) >= 11'sh0 & $signed(inSpriteYPreScaled_62) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1674 = {{1{inSpriteYPreScaled_62[10]}},inSpriteYPreScaled_62}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_63 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_63); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_63 = $signed(inSpriteXValue_63) >= 12'sh0 & $signed(inSpriteXValue_63) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1682 = {{1{inSpriteXValue_63[11]}},inSpriteXValue_63}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1877 = {{1{spriteYPositionReg_63[9]}},spriteYPositionReg_63}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_63 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1877); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_63 = inSpriteYValue_63[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_63 = $signed(inSpriteYPreScaled_63) >= 11'sh0 & $signed(inSpriteYPreScaled_63) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1690 = {{1{inSpriteYPreScaled_63[10]}},inSpriteYPreScaled_63}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteX_0 = _GEN_674[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_0 = _GEN_682[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_0_io_address_T_2 = 6'h20 * inSpriteY_0[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1881 = {{6'd0}, inSpriteX_0[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_0_io_address_T_4 = _GEN_1881 + _spriteMemories_0_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_3 = _GEN_722[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_3 = _GEN_730[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_3_io_address_T_2 = 6'h20 * inSpriteY_3[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1890 = {{6'd0}, inSpriteX_3[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_3_io_address_T_4 = _GEN_1890 + _spriteMemories_3_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_7 = _GEN_786[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_7 = _GEN_794[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_7_io_address_T_2 = 6'h20 * inSpriteY_7[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1902 = {{6'd0}, inSpriteX_7[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_7_io_address_T_4 = _GEN_1902 + _spriteMemories_7_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_8 = _GEN_802[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_8 = _GEN_810[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_8_io_address_T_2 = 6'h20 * inSpriteY_8[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1905 = {{6'd0}, inSpriteX_8[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_8_io_address_T_4 = _GEN_1905 + _spriteMemories_8_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_9 = _GEN_818[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_9 = _GEN_826[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_9_io_address_T_2 = 6'h20 * inSpriteY_9[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1908 = {{6'd0}, inSpriteX_9[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_9_io_address_T_4 = _GEN_1908 + _spriteMemories_9_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_10 = _GEN_834[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_10 = _GEN_842[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_10_io_address_T_2 = 6'h20 * inSpriteY_10[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1911 = {{6'd0}, inSpriteX_10[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_10_io_address_T_4 = _GEN_1911 + _spriteMemories_10_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_11 = _GEN_850[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_11 = _GEN_858[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_11_io_address_T_2 = 6'h20 * inSpriteY_11[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1914 = {{6'd0}, inSpriteX_11[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_11_io_address_T_4 = _GEN_1914 + _spriteMemories_11_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_12 = _GEN_866[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_12 = _GEN_874[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_12_io_address_T_2 = 6'h20 * inSpriteY_12[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1917 = {{6'd0}, inSpriteX_12[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_12_io_address_T_4 = _GEN_1917 + _spriteMemories_12_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_13 = _GEN_882[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_13 = _GEN_890[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_13_io_address_T_2 = 6'h20 * inSpriteY_13[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1920 = {{6'd0}, inSpriteX_13[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_13_io_address_T_4 = _GEN_1920 + _spriteMemories_13_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_14 = _GEN_898[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_14 = _GEN_906[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_14_io_address_T_2 = 6'h20 * inSpriteY_14[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1923 = {{6'd0}, inSpriteX_14[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_14_io_address_T_4 = _GEN_1923 + _spriteMemories_14_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_16 = _GEN_930[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_16 = _GEN_938[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_16_io_address_T_2 = 6'h20 * inSpriteY_16[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1929 = {{6'd0}, inSpriteX_16[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_16_io_address_T_4 = _GEN_1929 + _spriteMemories_16_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_17 = _GEN_946[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_17 = _GEN_954[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_17_io_address_T_2 = 6'h20 * inSpriteY_17[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1932 = {{6'd0}, inSpriteX_17[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_17_io_address_T_4 = _GEN_1932 + _spriteMemories_17_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_18 = _GEN_962[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_18 = _GEN_970[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_18_io_address_T_2 = 6'h20 * inSpriteY_18[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1935 = {{6'd0}, inSpriteX_18[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_18_io_address_T_4 = _GEN_1935 + _spriteMemories_18_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_19 = _GEN_978[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_19 = _GEN_986[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_19_io_address_T_2 = 6'h20 * inSpriteY_19[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1938 = {{6'd0}, inSpriteX_19[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_19_io_address_T_4 = _GEN_1938 + _spriteMemories_19_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_20 = _GEN_994[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_20 = _GEN_1002[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_20_io_address_T_2 = 6'h20 * inSpriteY_20[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1941 = {{6'd0}, inSpriteX_20[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_20_io_address_T_4 = _GEN_1941 + _spriteMemories_20_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_21 = _GEN_1010[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_21 = _GEN_1018[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_21_io_address_T_2 = 6'h20 * inSpriteY_21[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1944 = {{6'd0}, inSpriteX_21[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_21_io_address_T_4 = _GEN_1944 + _spriteMemories_21_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_22 = _GEN_1026[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_22 = _GEN_1034[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_22_io_address_T_2 = 6'h20 * inSpriteY_22[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1947 = {{6'd0}, inSpriteX_22[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_22_io_address_T_4 = _GEN_1947 + _spriteMemories_22_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_23 = _GEN_1042[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_23 = _GEN_1050[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_23_io_address_T_2 = 6'h20 * inSpriteY_23[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1950 = {{6'd0}, inSpriteX_23[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_23_io_address_T_4 = _GEN_1950 + _spriteMemories_23_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_24 = _GEN_1058[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_24 = _GEN_1066[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_24_io_address_T_2 = 6'h20 * inSpriteY_24[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1953 = {{6'd0}, inSpriteX_24[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_24_io_address_T_4 = _GEN_1953 + _spriteMemories_24_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_25 = _GEN_1074[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_25 = _GEN_1082[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_25_io_address_T_2 = 6'h20 * inSpriteY_25[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1956 = {{6'd0}, inSpriteX_25[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_25_io_address_T_4 = _GEN_1956 + _spriteMemories_25_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_26 = _GEN_1090[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_26 = _GEN_1098[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_26_io_address_T_2 = 6'h20 * inSpriteY_26[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1959 = {{6'd0}, inSpriteX_26[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_26_io_address_T_4 = _GEN_1959 + _spriteMemories_26_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_27 = _GEN_1106[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_27 = _GEN_1114[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_27_io_address_T_2 = 6'h20 * inSpriteY_27[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1962 = {{6'd0}, inSpriteX_27[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_27_io_address_T_4 = _GEN_1962 + _spriteMemories_27_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_28 = _GEN_1122[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_28 = _GEN_1130[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_28_io_address_T_2 = 6'h20 * inSpriteY_28[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1965 = {{6'd0}, inSpriteX_28[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_28_io_address_T_4 = _GEN_1965 + _spriteMemories_28_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_29 = _GEN_1138[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_29 = _GEN_1146[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_29_io_address_T_2 = 6'h20 * inSpriteY_29[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1968 = {{6'd0}, inSpriteX_29[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_29_io_address_T_4 = _GEN_1968 + _spriteMemories_29_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_30 = _GEN_1154[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_30 = _GEN_1162[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_30_io_address_T_2 = 6'h20 * inSpriteY_30[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1971 = {{6'd0}, inSpriteX_30[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_30_io_address_T_4 = _GEN_1971 + _spriteMemories_30_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_31 = _GEN_1170[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_31 = _GEN_1178[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_31_io_address_T_2 = 6'h20 * inSpriteY_31[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1974 = {{6'd0}, inSpriteX_31[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_31_io_address_T_4 = _GEN_1974 + _spriteMemories_31_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_32 = _GEN_1186[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_32 = _GEN_1194[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_32_io_address_T_2 = 6'h20 * inSpriteY_32[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1977 = {{6'd0}, inSpriteX_32[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_32_io_address_T_4 = _GEN_1977 + _spriteMemories_32_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_33 = _GEN_1202[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_33 = _GEN_1210[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_33_io_address_T_2 = 6'h20 * inSpriteY_33[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1980 = {{6'd0}, inSpriteX_33[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_33_io_address_T_4 = _GEN_1980 + _spriteMemories_33_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_34 = _GEN_1218[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_34 = _GEN_1226[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_34_io_address_T_2 = 6'h20 * inSpriteY_34[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1983 = {{6'd0}, inSpriteX_34[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_34_io_address_T_4 = _GEN_1983 + _spriteMemories_34_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_35 = _GEN_1234[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_35 = _GEN_1242[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_35_io_address_T_2 = 6'h20 * inSpriteY_35[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1986 = {{6'd0}, inSpriteX_35[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_35_io_address_T_4 = _GEN_1986 + _spriteMemories_35_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_36 = _GEN_1250[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_36 = _GEN_1258[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_36_io_address_T_2 = 6'h20 * inSpriteY_36[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1989 = {{6'd0}, inSpriteX_36[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_36_io_address_T_4 = _GEN_1989 + _spriteMemories_36_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_37 = _GEN_1266[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_37 = _GEN_1274[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_37_io_address_T_2 = 6'h20 * inSpriteY_37[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1992 = {{6'd0}, inSpriteX_37[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_37_io_address_T_4 = _GEN_1992 + _spriteMemories_37_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_38 = _GEN_1282[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_38 = _GEN_1290[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_38_io_address_T_2 = 6'h20 * inSpriteY_38[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1995 = {{6'd0}, inSpriteX_38[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_38_io_address_T_4 = _GEN_1995 + _spriteMemories_38_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_39 = _GEN_1298[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_39 = _GEN_1306[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_39_io_address_T_2 = 6'h20 * inSpriteY_39[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1998 = {{6'd0}, inSpriteX_39[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_39_io_address_T_4 = _GEN_1998 + _spriteMemories_39_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_40 = _GEN_1314[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_40 = _GEN_1322[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_40_io_address_T_2 = 6'h20 * inSpriteY_40[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2001 = {{6'd0}, inSpriteX_40[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_40_io_address_T_4 = _GEN_2001 + _spriteMemories_40_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_41 = _GEN_1330[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_41 = _GEN_1338[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_41_io_address_T_2 = 6'h20 * inSpriteY_41[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2004 = {{6'd0}, inSpriteX_41[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_41_io_address_T_4 = _GEN_2004 + _spriteMemories_41_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_42 = _GEN_1346[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_42 = _GEN_1354[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_42_io_address_T_2 = 6'h20 * inSpriteY_42[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2007 = {{6'd0}, inSpriteX_42[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_42_io_address_T_4 = _GEN_2007 + _spriteMemories_42_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_43 = _GEN_1362[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_43 = _GEN_1370[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_43_io_address_T_2 = 6'h20 * inSpriteY_43[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2010 = {{6'd0}, inSpriteX_43[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_43_io_address_T_4 = _GEN_2010 + _spriteMemories_43_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_44 = _GEN_1378[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_44 = _GEN_1386[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_44_io_address_T_2 = 6'h20 * inSpriteY_44[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2013 = {{6'd0}, inSpriteX_44[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_44_io_address_T_4 = _GEN_2013 + _spriteMemories_44_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_45 = _GEN_1394[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_45 = _GEN_1402[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_45_io_address_T_2 = 6'h20 * inSpriteY_45[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2016 = {{6'd0}, inSpriteX_45[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_45_io_address_T_4 = _GEN_2016 + _spriteMemories_45_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_46 = _GEN_1410[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_46 = _GEN_1418[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_46_io_address_T_2 = 6'h20 * inSpriteY_46[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2019 = {{6'd0}, inSpriteX_46[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_46_io_address_T_4 = _GEN_2019 + _spriteMemories_46_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_47 = _GEN_1426[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_47 = _GEN_1434[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_47_io_address_T_2 = 6'h20 * inSpriteY_47[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2022 = {{6'd0}, inSpriteX_47[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_47_io_address_T_4 = _GEN_2022 + _spriteMemories_47_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_48 = _GEN_1442[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_48 = _GEN_1450[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_48_io_address_T_2 = 6'h20 * inSpriteY_48[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2025 = {{6'd0}, inSpriteX_48[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_48_io_address_T_4 = _GEN_2025 + _spriteMemories_48_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_49 = _GEN_1458[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_49 = _GEN_1466[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_49_io_address_T_2 = 6'h20 * inSpriteY_49[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2028 = {{6'd0}, inSpriteX_49[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_49_io_address_T_4 = _GEN_2028 + _spriteMemories_49_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_50 = _GEN_1474[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_50 = _GEN_1482[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_50_io_address_T_2 = 6'h20 * inSpriteY_50[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2031 = {{6'd0}, inSpriteX_50[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_50_io_address_T_4 = _GEN_2031 + _spriteMemories_50_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_51 = _GEN_1490[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_51 = _GEN_1498[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_51_io_address_T_2 = 6'h20 * inSpriteY_51[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2034 = {{6'd0}, inSpriteX_51[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_51_io_address_T_4 = _GEN_2034 + _spriteMemories_51_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_52 = _GEN_1506[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_52 = _GEN_1514[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_52_io_address_T_2 = 6'h20 * inSpriteY_52[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2037 = {{6'd0}, inSpriteX_52[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_52_io_address_T_4 = _GEN_2037 + _spriteMemories_52_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_53 = _GEN_1522[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_53 = _GEN_1530[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_53_io_address_T_2 = 6'h20 * inSpriteY_53[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2040 = {{6'd0}, inSpriteX_53[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_53_io_address_T_4 = _GEN_2040 + _spriteMemories_53_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_54 = _GEN_1538[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_54 = _GEN_1546[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_54_io_address_T_2 = 6'h20 * inSpriteY_54[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2043 = {{6'd0}, inSpriteX_54[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_54_io_address_T_4 = _GEN_2043 + _spriteMemories_54_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_55 = _GEN_1554[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_55 = _GEN_1562[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_55_io_address_T_2 = 6'h20 * inSpriteY_55[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2046 = {{6'd0}, inSpriteX_55[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_55_io_address_T_4 = _GEN_2046 + _spriteMemories_55_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_56 = _GEN_1570[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_56 = _GEN_1578[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_56_io_address_T_2 = 6'h20 * inSpriteY_56[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2049 = {{6'd0}, inSpriteX_56[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_56_io_address_T_4 = _GEN_2049 + _spriteMemories_56_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_57 = _GEN_1586[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_57 = _GEN_1594[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_57_io_address_T_2 = 6'h20 * inSpriteY_57[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2052 = {{6'd0}, inSpriteX_57[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_57_io_address_T_4 = _GEN_2052 + _spriteMemories_57_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_58 = _GEN_1602[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_58 = _GEN_1610[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_58_io_address_T_2 = 6'h20 * inSpriteY_58[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2055 = {{6'd0}, inSpriteX_58[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_58_io_address_T_4 = _GEN_2055 + _spriteMemories_58_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_59 = _GEN_1618[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_59 = _GEN_1626[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_59_io_address_T_2 = 6'h20 * inSpriteY_59[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2058 = {{6'd0}, inSpriteX_59[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_59_io_address_T_4 = _GEN_2058 + _spriteMemories_59_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_60 = _GEN_1634[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_60 = _GEN_1642[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_60_io_address_T_2 = 6'h20 * inSpriteY_60[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2061 = {{6'd0}, inSpriteX_60[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_60_io_address_T_4 = _GEN_2061 + _spriteMemories_60_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_61 = _GEN_1650[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_61 = _GEN_1658[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_61_io_address_T_2 = 6'h20 * inSpriteY_61[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2064 = {{6'd0}, inSpriteX_61[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_61_io_address_T_4 = _GEN_2064 + _spriteMemories_61_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_62 = _GEN_1666[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_62 = _GEN_1674[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_62_io_address_T_2 = 6'h20 * inSpriteY_62[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2067 = {{6'd0}, inSpriteX_62[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_62_io_address_T_4 = _GEN_2067 + _spriteMemories_62_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_63 = _GEN_1682[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_63 = _GEN_1690[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_63_io_address_T_2 = 6'h20 * inSpriteY_63[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2070 = {{6'd0}, inSpriteX_63[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_63_io_address_T_4 = _GEN_2070 + _spriteMemories_63_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] pixelColorSprite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 339:33]
  reg  pixelColorSpriteValid; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 340:38]
  wire [5:0] pixelColorInDisplay = pixelColorSpriteValid ? pixelColorSprite : pixelColorBack; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 344:32]
  reg  pixelColourVGA_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  pixelColourVGA_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  pixelColourVGA_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  wire [5:0] pixelColourVGA = pixelColourVGA_pipeReg_0 ? pixelColorInDisplay : 6'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 345:27]
  reg [3:0] io_vgaRed_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 349:23]
  reg [3:0] io_vgaGreen_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 350:25]
  reg [3:0] io_vgaBlue_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 351:24]
  Memory backTileMemories_0 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_0_clock),
    .io_address(backTileMemories_0_io_address),
    .io_dataRead(backTileMemories_0_io_dataRead)
  );
  Memory_1 backTileMemories_1 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_1_clock),
    .io_address(backTileMemories_1_io_address),
    .io_dataRead(backTileMemories_1_io_dataRead)
  );
  Memory_2 backTileMemories_2 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_2_clock),
    .io_address(backTileMemories_2_io_address),
    .io_dataRead(backTileMemories_2_io_dataRead)
  );
  Memory_3 backTileMemories_3 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_3_clock),
    .io_address(backTileMemories_3_io_address),
    .io_dataRead(backTileMemories_3_io_dataRead)
  );
  Memory_4 backTileMemories_4 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_4_clock),
    .io_address(backTileMemories_4_io_address),
    .io_dataRead(backTileMemories_4_io_dataRead)
  );
  Memory_5 backTileMemories_5 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_5_clock),
    .io_address(backTileMemories_5_io_address),
    .io_dataRead(backTileMemories_5_io_dataRead)
  );
  Memory_6 backTileMemories_6 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_6_clock),
    .io_address(backTileMemories_6_io_address),
    .io_dataRead(backTileMemories_6_io_dataRead)
  );
  Memory_7 backTileMemories_7 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_7_clock),
    .io_address(backTileMemories_7_io_address),
    .io_dataRead(backTileMemories_7_io_dataRead)
  );
  Memory_8 backTileMemories_8 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_8_clock),
    .io_address(backTileMemories_8_io_address),
    .io_dataRead(backTileMemories_8_io_dataRead)
  );
  Memory_9 backTileMemories_9 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_9_clock),
    .io_address(backTileMemories_9_io_address),
    .io_dataRead(backTileMemories_9_io_dataRead)
  );
  Memory_10 backTileMemories_10 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_10_clock),
    .io_address(backTileMemories_10_io_address),
    .io_dataRead(backTileMemories_10_io_dataRead)
  );
  Memory_11 backTileMemories_11 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_11_clock),
    .io_address(backTileMemories_11_io_address),
    .io_dataRead(backTileMemories_11_io_dataRead)
  );
  Memory_12 backTileMemories_12 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_12_clock),
    .io_address(backTileMemories_12_io_address),
    .io_dataRead(backTileMemories_12_io_dataRead)
  );
  Memory_13 backTileMemories_13 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_13_clock),
    .io_address(backTileMemories_13_io_address),
    .io_dataRead(backTileMemories_13_io_dataRead)
  );
  Memory_14 backTileMemories_14 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_14_clock),
    .io_address(backTileMemories_14_io_address),
    .io_dataRead(backTileMemories_14_io_dataRead)
  );
  Memory_15 backTileMemories_15 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_15_clock),
    .io_address(backTileMemories_15_io_address),
    .io_dataRead(backTileMemories_15_io_dataRead)
  );
  Memory_16 backTileMemories_16 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_16_clock),
    .io_address(backTileMemories_16_io_address),
    .io_dataRead(backTileMemories_16_io_dataRead)
  );
  Memory_17 backTileMemories_17 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_17_clock),
    .io_address(backTileMemories_17_io_address),
    .io_dataRead(backTileMemories_17_io_dataRead)
  );
  Memory_18 backTileMemories_18 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_18_clock),
    .io_address(backTileMemories_18_io_address),
    .io_dataRead(backTileMemories_18_io_dataRead)
  );
  Memory_19 backTileMemories_19 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_19_clock),
    .io_address(backTileMemories_19_io_address),
    .io_dataRead(backTileMemories_19_io_dataRead)
  );
  Memory_20 backTileMemories_20 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_20_clock),
    .io_address(backTileMemories_20_io_address),
    .io_dataRead(backTileMemories_20_io_dataRead)
  );
  Memory_21 backTileMemories_21 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_21_clock),
    .io_address(backTileMemories_21_io_address),
    .io_dataRead(backTileMemories_21_io_dataRead)
  );
  Memory_22 backTileMemories_22 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_22_clock),
    .io_address(backTileMemories_22_io_address),
    .io_dataRead(backTileMemories_22_io_dataRead)
  );
  Memory_23 backTileMemories_23 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_23_clock),
    .io_address(backTileMemories_23_io_address),
    .io_dataRead(backTileMemories_23_io_dataRead)
  );
  Memory_24 backTileMemories_24 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_24_clock),
    .io_address(backTileMemories_24_io_address),
    .io_dataRead(backTileMemories_24_io_dataRead)
  );
  Memory_25 backTileMemories_25 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_25_clock),
    .io_address(backTileMemories_25_io_address),
    .io_dataRead(backTileMemories_25_io_dataRead)
  );
  Memory_26 backTileMemories_26 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_26_clock),
    .io_address(backTileMemories_26_io_address),
    .io_dataRead(backTileMemories_26_io_dataRead)
  );
  Memory_27 backTileMemories_27 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_27_clock),
    .io_address(backTileMemories_27_io_address),
    .io_dataRead(backTileMemories_27_io_dataRead)
  );
  Memory_28 backTileMemories_28 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_28_clock),
    .io_address(backTileMemories_28_io_address),
    .io_dataRead(backTileMemories_28_io_dataRead)
  );
  Memory_29 backTileMemories_29 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_29_clock),
    .io_address(backTileMemories_29_io_address),
    .io_dataRead(backTileMemories_29_io_dataRead)
  );
  Memory_30 backTileMemories_30 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_30_clock),
    .io_address(backTileMemories_30_io_address),
    .io_dataRead(backTileMemories_30_io_dataRead)
  );
  Memory_31 backTileMemories_31 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_31_clock),
    .io_address(backTileMemories_31_io_address),
    .io_dataRead(backTileMemories_31_io_dataRead)
  );
  Memory_32 backTileMemories_32 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_32_clock),
    .io_address(backTileMemories_32_io_address),
    .io_dataRead(backTileMemories_32_io_dataRead)
  );
  Memory_33 backTileMemories_33 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_33_clock),
    .io_address(backTileMemories_33_io_address),
    .io_dataRead(backTileMemories_33_io_dataRead)
  );
  Memory_34 backTileMemories_34 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_34_clock),
    .io_address(backTileMemories_34_io_address),
    .io_dataRead(backTileMemories_34_io_dataRead)
  );
  Memory_35 backTileMemories_35 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_35_clock),
    .io_address(backTileMemories_35_io_address),
    .io_dataRead(backTileMemories_35_io_dataRead)
  );
  Memory_36 backTileMemories_36 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_36_clock),
    .io_address(backTileMemories_36_io_address),
    .io_dataRead(backTileMemories_36_io_dataRead)
  );
  Memory_37 backTileMemories_37 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_37_clock),
    .io_address(backTileMemories_37_io_address),
    .io_dataRead(backTileMemories_37_io_dataRead)
  );
  Memory_38 backTileMemories_38 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_38_clock),
    .io_address(backTileMemories_38_io_address),
    .io_dataRead(backTileMemories_38_io_dataRead)
  );
  Memory_39 backTileMemories_39 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_39_clock),
    .io_address(backTileMemories_39_io_address),
    .io_dataRead(backTileMemories_39_io_dataRead)
  );
  Memory_40 backTileMemories_40 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_40_clock),
    .io_address(backTileMemories_40_io_address),
    .io_dataRead(backTileMemories_40_io_dataRead)
  );
  Memory_41 backTileMemories_41 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_41_clock),
    .io_address(backTileMemories_41_io_address),
    .io_dataRead(backTileMemories_41_io_dataRead)
  );
  Memory_42 backTileMemories_42 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_42_clock),
    .io_address(backTileMemories_42_io_address),
    .io_dataRead(backTileMemories_42_io_dataRead)
  );
  Memory_43 backTileMemories_43 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_43_clock),
    .io_address(backTileMemories_43_io_address),
    .io_dataRead(backTileMemories_43_io_dataRead)
  );
  Memory_44 backTileMemories_44 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_44_clock),
    .io_address(backTileMemories_44_io_address),
    .io_dataRead(backTileMemories_44_io_dataRead)
  );
  Memory_45 backTileMemories_45 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_45_clock),
    .io_address(backTileMemories_45_io_address),
    .io_dataRead(backTileMemories_45_io_dataRead)
  );
  Memory_46 backTileMemories_46 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_46_clock),
    .io_address(backTileMemories_46_io_address),
    .io_dataRead(backTileMemories_46_io_dataRead)
  );
  Memory_47 backTileMemories_47 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_47_clock),
    .io_address(backTileMemories_47_io_address),
    .io_dataRead(backTileMemories_47_io_dataRead)
  );
  Memory_48 backTileMemories_48 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_48_clock),
    .io_address(backTileMemories_48_io_address),
    .io_dataRead(backTileMemories_48_io_dataRead)
  );
  Memory_49 backTileMemories_49 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_49_clock),
    .io_address(backTileMemories_49_io_address),
    .io_dataRead(backTileMemories_49_io_dataRead)
  );
  Memory_50 backTileMemories_50 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_50_clock),
    .io_address(backTileMemories_50_io_address),
    .io_dataRead(backTileMemories_50_io_dataRead)
  );
  Memory_51 backTileMemories_51 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_51_clock),
    .io_address(backTileMemories_51_io_address),
    .io_dataRead(backTileMemories_51_io_dataRead)
  );
  Memory_52 backTileMemories_52 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_52_clock),
    .io_address(backTileMemories_52_io_address),
    .io_dataRead(backTileMemories_52_io_dataRead)
  );
  Memory_53 backTileMemories_53 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_53_clock),
    .io_address(backTileMemories_53_io_address),
    .io_dataRead(backTileMemories_53_io_dataRead)
  );
  Memory_54 backTileMemories_54 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_54_clock),
    .io_address(backTileMemories_54_io_address),
    .io_dataRead(backTileMemories_54_io_dataRead)
  );
  Memory_55 backTileMemories_55 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_55_clock),
    .io_address(backTileMemories_55_io_address),
    .io_dataRead(backTileMemories_55_io_dataRead)
  );
  Memory_56 backTileMemories_56 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_56_clock),
    .io_address(backTileMemories_56_io_address),
    .io_dataRead(backTileMemories_56_io_dataRead)
  );
  Memory_57 backTileMemories_57 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_57_clock),
    .io_address(backTileMemories_57_io_address),
    .io_dataRead(backTileMemories_57_io_dataRead)
  );
  Memory_58 backTileMemories_58 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_58_clock),
    .io_address(backTileMemories_58_io_address),
    .io_dataRead(backTileMemories_58_io_dataRead)
  );
  Memory_59 backTileMemories_59 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_59_clock),
    .io_address(backTileMemories_59_io_address),
    .io_dataRead(backTileMemories_59_io_dataRead)
  );
  Memory_60 backTileMemories_60 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_60_clock),
    .io_address(backTileMemories_60_io_address),
    .io_dataRead(backTileMemories_60_io_dataRead)
  );
  Memory_61 backTileMemories_61 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_61_clock),
    .io_address(backTileMemories_61_io_address),
    .io_dataRead(backTileMemories_61_io_dataRead)
  );
  Memory_62 backTileMemories_62 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_62_clock),
    .io_address(backTileMemories_62_io_address),
    .io_dataRead(backTileMemories_62_io_dataRead)
  );
  Memory_63 backTileMemories_63 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_63_clock),
    .io_address(backTileMemories_63_io_address),
    .io_dataRead(backTileMemories_63_io_dataRead)
  );
  Memory_64 backBufferMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
    .clock(backBufferMemory_clock),
    .io_address(backBufferMemory_io_address),
    .io_dataRead(backBufferMemory_io_dataRead),
    .io_writeEnable(backBufferMemory_io_writeEnable),
    .io_dataWrite(backBufferMemory_io_dataWrite)
  );
  Memory_64 backBufferShadowMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
    .clock(backBufferShadowMemory_clock),
    .io_address(backBufferShadowMemory_io_address),
    .io_dataRead(backBufferShadowMemory_io_dataRead),
    .io_writeEnable(backBufferShadowMemory_io_writeEnable),
    .io_dataWrite(backBufferShadowMemory_io_dataWrite)
  );
  Memory_66 backBufferRestoreMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
    .clock(backBufferRestoreMemory_clock),
    .io_address(backBufferRestoreMemory_io_address),
    .io_dataRead(backBufferRestoreMemory_io_dataRead)
  );
  Memory_67 spriteMemories_0 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_0_clock),
    .io_address(spriteMemories_0_io_address),
    .io_dataRead(spriteMemories_0_io_dataRead)
  );
  Memory_68 spriteMemories_1 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_1_clock),
    .io_address(spriteMemories_1_io_address),
    .io_dataRead(spriteMemories_1_io_dataRead)
  );
  Memory_69 spriteMemories_2 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_2_clock),
    .io_address(spriteMemories_2_io_address),
    .io_dataRead(spriteMemories_2_io_dataRead)
  );
  Memory_70 spriteMemories_3 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_3_clock),
    .io_address(spriteMemories_3_io_address),
    .io_dataRead(spriteMemories_3_io_dataRead)
  );
  Memory_71 spriteMemories_4 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_4_clock),
    .io_address(spriteMemories_4_io_address),
    .io_dataRead(spriteMemories_4_io_dataRead)
  );
  Memory_72 spriteMemories_5 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_5_clock),
    .io_address(spriteMemories_5_io_address),
    .io_dataRead(spriteMemories_5_io_dataRead)
  );
  Memory_73 spriteMemories_6 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_6_clock),
    .io_address(spriteMemories_6_io_address),
    .io_dataRead(spriteMemories_6_io_dataRead)
  );
  Memory_74 spriteMemories_7 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_7_clock),
    .io_address(spriteMemories_7_io_address),
    .io_dataRead(spriteMemories_7_io_dataRead)
  );
  Memory_75 spriteMemories_8 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_8_clock),
    .io_address(spriteMemories_8_io_address),
    .io_dataRead(spriteMemories_8_io_dataRead)
  );
  Memory_76 spriteMemories_9 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_9_clock),
    .io_address(spriteMemories_9_io_address),
    .io_dataRead(spriteMemories_9_io_dataRead)
  );
  Memory_77 spriteMemories_10 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_10_clock),
    .io_address(spriteMemories_10_io_address),
    .io_dataRead(spriteMemories_10_io_dataRead)
  );
  Memory_78 spriteMemories_11 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_11_clock),
    .io_address(spriteMemories_11_io_address),
    .io_dataRead(spriteMemories_11_io_dataRead)
  );
  Memory_79 spriteMemories_12 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_12_clock),
    .io_address(spriteMemories_12_io_address),
    .io_dataRead(spriteMemories_12_io_dataRead)
  );
  Memory_80 spriteMemories_13 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_13_clock),
    .io_address(spriteMemories_13_io_address),
    .io_dataRead(spriteMemories_13_io_dataRead)
  );
  Memory_81 spriteMemories_14 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_14_clock),
    .io_address(spriteMemories_14_io_address),
    .io_dataRead(spriteMemories_14_io_dataRead)
  );
  Memory_82 spriteMemories_15 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_15_clock),
    .io_address(spriteMemories_15_io_address),
    .io_dataRead(spriteMemories_15_io_dataRead)
  );
  Memory_83 spriteMemories_16 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_16_clock),
    .io_address(spriteMemories_16_io_address),
    .io_dataRead(spriteMemories_16_io_dataRead)
  );
  Memory_84 spriteMemories_17 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_17_clock),
    .io_address(spriteMemories_17_io_address),
    .io_dataRead(spriteMemories_17_io_dataRead)
  );
  Memory_85 spriteMemories_18 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_18_clock),
    .io_address(spriteMemories_18_io_address),
    .io_dataRead(spriteMemories_18_io_dataRead)
  );
  Memory_86 spriteMemories_19 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_19_clock),
    .io_address(spriteMemories_19_io_address),
    .io_dataRead(spriteMemories_19_io_dataRead)
  );
  Memory_87 spriteMemories_20 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_20_clock),
    .io_address(spriteMemories_20_io_address),
    .io_dataRead(spriteMemories_20_io_dataRead)
  );
  Memory_88 spriteMemories_21 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_21_clock),
    .io_address(spriteMemories_21_io_address),
    .io_dataRead(spriteMemories_21_io_dataRead)
  );
  Memory_89 spriteMemories_22 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_22_clock),
    .io_address(spriteMemories_22_io_address),
    .io_dataRead(spriteMemories_22_io_dataRead)
  );
  Memory_90 spriteMemories_23 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_23_clock),
    .io_address(spriteMemories_23_io_address),
    .io_dataRead(spriteMemories_23_io_dataRead)
  );
  Memory_91 spriteMemories_24 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_24_clock),
    .io_address(spriteMemories_24_io_address),
    .io_dataRead(spriteMemories_24_io_dataRead)
  );
  Memory_92 spriteMemories_25 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_25_clock),
    .io_address(spriteMemories_25_io_address),
    .io_dataRead(spriteMemories_25_io_dataRead)
  );
  Memory_93 spriteMemories_26 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_26_clock),
    .io_address(spriteMemories_26_io_address),
    .io_dataRead(spriteMemories_26_io_dataRead)
  );
  Memory_94 spriteMemories_27 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_27_clock),
    .io_address(spriteMemories_27_io_address),
    .io_dataRead(spriteMemories_27_io_dataRead)
  );
  Memory_95 spriteMemories_28 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_28_clock),
    .io_address(spriteMemories_28_io_address),
    .io_dataRead(spriteMemories_28_io_dataRead)
  );
  Memory_96 spriteMemories_29 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_29_clock),
    .io_address(spriteMemories_29_io_address),
    .io_dataRead(spriteMemories_29_io_dataRead)
  );
  Memory_97 spriteMemories_30 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_30_clock),
    .io_address(spriteMemories_30_io_address),
    .io_dataRead(spriteMemories_30_io_dataRead)
  );
  Memory_98 spriteMemories_31 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_31_clock),
    .io_address(spriteMemories_31_io_address),
    .io_dataRead(spriteMemories_31_io_dataRead)
  );
  Memory_99 spriteMemories_32 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_32_clock),
    .io_address(spriteMemories_32_io_address),
    .io_dataRead(spriteMemories_32_io_dataRead)
  );
  Memory_100 spriteMemories_33 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_33_clock),
    .io_address(spriteMemories_33_io_address),
    .io_dataRead(spriteMemories_33_io_dataRead)
  );
  Memory_101 spriteMemories_34 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_34_clock),
    .io_address(spriteMemories_34_io_address),
    .io_dataRead(spriteMemories_34_io_dataRead)
  );
  Memory_102 spriteMemories_35 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_35_clock),
    .io_address(spriteMemories_35_io_address),
    .io_dataRead(spriteMemories_35_io_dataRead)
  );
  Memory_103 spriteMemories_36 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_36_clock),
    .io_address(spriteMemories_36_io_address),
    .io_dataRead(spriteMemories_36_io_dataRead)
  );
  Memory_104 spriteMemories_37 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_37_clock),
    .io_address(spriteMemories_37_io_address),
    .io_dataRead(spriteMemories_37_io_dataRead)
  );
  Memory_105 spriteMemories_38 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_38_clock),
    .io_address(spriteMemories_38_io_address),
    .io_dataRead(spriteMemories_38_io_dataRead)
  );
  Memory_106 spriteMemories_39 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_39_clock),
    .io_address(spriteMemories_39_io_address),
    .io_dataRead(spriteMemories_39_io_dataRead)
  );
  Memory_107 spriteMemories_40 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_40_clock),
    .io_address(spriteMemories_40_io_address),
    .io_dataRead(spriteMemories_40_io_dataRead)
  );
  Memory_108 spriteMemories_41 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_41_clock),
    .io_address(spriteMemories_41_io_address),
    .io_dataRead(spriteMemories_41_io_dataRead)
  );
  Memory_109 spriteMemories_42 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_42_clock),
    .io_address(spriteMemories_42_io_address),
    .io_dataRead(spriteMemories_42_io_dataRead)
  );
  Memory_110 spriteMemories_43 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_43_clock),
    .io_address(spriteMemories_43_io_address),
    .io_dataRead(spriteMemories_43_io_dataRead)
  );
  Memory_111 spriteMemories_44 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_44_clock),
    .io_address(spriteMemories_44_io_address),
    .io_dataRead(spriteMemories_44_io_dataRead)
  );
  Memory_112 spriteMemories_45 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_45_clock),
    .io_address(spriteMemories_45_io_address),
    .io_dataRead(spriteMemories_45_io_dataRead)
  );
  Memory_113 spriteMemories_46 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_46_clock),
    .io_address(spriteMemories_46_io_address),
    .io_dataRead(spriteMemories_46_io_dataRead)
  );
  Memory_114 spriteMemories_47 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_47_clock),
    .io_address(spriteMemories_47_io_address),
    .io_dataRead(spriteMemories_47_io_dataRead)
  );
  Memory_115 spriteMemories_48 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_48_clock),
    .io_address(spriteMemories_48_io_address),
    .io_dataRead(spriteMemories_48_io_dataRead)
  );
  Memory_116 spriteMemories_49 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_49_clock),
    .io_address(spriteMemories_49_io_address),
    .io_dataRead(spriteMemories_49_io_dataRead)
  );
  Memory_117 spriteMemories_50 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_50_clock),
    .io_address(spriteMemories_50_io_address),
    .io_dataRead(spriteMemories_50_io_dataRead)
  );
  Memory_118 spriteMemories_51 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_51_clock),
    .io_address(spriteMemories_51_io_address),
    .io_dataRead(spriteMemories_51_io_dataRead)
  );
  Memory_119 spriteMemories_52 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_52_clock),
    .io_address(spriteMemories_52_io_address),
    .io_dataRead(spriteMemories_52_io_dataRead)
  );
  Memory_120 spriteMemories_53 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_53_clock),
    .io_address(spriteMemories_53_io_address),
    .io_dataRead(spriteMemories_53_io_dataRead)
  );
  Memory_121 spriteMemories_54 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_54_clock),
    .io_address(spriteMemories_54_io_address),
    .io_dataRead(spriteMemories_54_io_dataRead)
  );
  Memory_122 spriteMemories_55 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_55_clock),
    .io_address(spriteMemories_55_io_address),
    .io_dataRead(spriteMemories_55_io_dataRead)
  );
  Memory_123 spriteMemories_56 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_56_clock),
    .io_address(spriteMemories_56_io_address),
    .io_dataRead(spriteMemories_56_io_dataRead)
  );
  Memory_124 spriteMemories_57 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_57_clock),
    .io_address(spriteMemories_57_io_address),
    .io_dataRead(spriteMemories_57_io_dataRead)
  );
  Memory_125 spriteMemories_58 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_58_clock),
    .io_address(spriteMemories_58_io_address),
    .io_dataRead(spriteMemories_58_io_dataRead)
  );
  Memory_126 spriteMemories_59 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_59_clock),
    .io_address(spriteMemories_59_io_address),
    .io_dataRead(spriteMemories_59_io_dataRead)
  );
  Memory_127 spriteMemories_60 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_60_clock),
    .io_address(spriteMemories_60_io_address),
    .io_dataRead(spriteMemories_60_io_dataRead)
  );
  Memory_128 spriteMemories_61 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_61_clock),
    .io_address(spriteMemories_61_io_address),
    .io_dataRead(spriteMemories_61_io_dataRead)
  );
  Memory_129 spriteMemories_62 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_62_clock),
    .io_address(spriteMemories_62_io_address),
    .io_dataRead(spriteMemories_62_io_dataRead)
  );
  Memory_130 spriteMemories_63 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_63_clock),
    .io_address(spriteMemories_63_io_address),
    .io_dataRead(spriteMemories_63_io_dataRead)
  );
  MultiHotPriortyReductionTree multiHotPriortyReductionTree ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
    .io_dataInput_0(multiHotPriortyReductionTree_io_dataInput_0),
    .io_dataInput_1(multiHotPriortyReductionTree_io_dataInput_1),
    .io_dataInput_2(multiHotPriortyReductionTree_io_dataInput_2),
    .io_dataInput_3(multiHotPriortyReductionTree_io_dataInput_3),
    .io_dataInput_4(multiHotPriortyReductionTree_io_dataInput_4),
    .io_dataInput_5(multiHotPriortyReductionTree_io_dataInput_5),
    .io_dataInput_6(multiHotPriortyReductionTree_io_dataInput_6),
    .io_dataInput_7(multiHotPriortyReductionTree_io_dataInput_7),
    .io_dataInput_8(multiHotPriortyReductionTree_io_dataInput_8),
    .io_dataInput_9(multiHotPriortyReductionTree_io_dataInput_9),
    .io_dataInput_10(multiHotPriortyReductionTree_io_dataInput_10),
    .io_dataInput_11(multiHotPriortyReductionTree_io_dataInput_11),
    .io_dataInput_12(multiHotPriortyReductionTree_io_dataInput_12),
    .io_dataInput_13(multiHotPriortyReductionTree_io_dataInput_13),
    .io_dataInput_14(multiHotPriortyReductionTree_io_dataInput_14),
    .io_dataInput_15(multiHotPriortyReductionTree_io_dataInput_15),
    .io_dataInput_16(multiHotPriortyReductionTree_io_dataInput_16),
    .io_dataInput_17(multiHotPriortyReductionTree_io_dataInput_17),
    .io_dataInput_18(multiHotPriortyReductionTree_io_dataInput_18),
    .io_dataInput_19(multiHotPriortyReductionTree_io_dataInput_19),
    .io_dataInput_20(multiHotPriortyReductionTree_io_dataInput_20),
    .io_dataInput_21(multiHotPriortyReductionTree_io_dataInput_21),
    .io_dataInput_22(multiHotPriortyReductionTree_io_dataInput_22),
    .io_dataInput_23(multiHotPriortyReductionTree_io_dataInput_23),
    .io_dataInput_24(multiHotPriortyReductionTree_io_dataInput_24),
    .io_dataInput_25(multiHotPriortyReductionTree_io_dataInput_25),
    .io_dataInput_26(multiHotPriortyReductionTree_io_dataInput_26),
    .io_dataInput_27(multiHotPriortyReductionTree_io_dataInput_27),
    .io_dataInput_28(multiHotPriortyReductionTree_io_dataInput_28),
    .io_dataInput_29(multiHotPriortyReductionTree_io_dataInput_29),
    .io_dataInput_30(multiHotPriortyReductionTree_io_dataInput_30),
    .io_dataInput_31(multiHotPriortyReductionTree_io_dataInput_31),
    .io_dataInput_32(multiHotPriortyReductionTree_io_dataInput_32),
    .io_dataInput_33(multiHotPriortyReductionTree_io_dataInput_33),
    .io_dataInput_34(multiHotPriortyReductionTree_io_dataInput_34),
    .io_dataInput_35(multiHotPriortyReductionTree_io_dataInput_35),
    .io_dataInput_36(multiHotPriortyReductionTree_io_dataInput_36),
    .io_dataInput_37(multiHotPriortyReductionTree_io_dataInput_37),
    .io_dataInput_38(multiHotPriortyReductionTree_io_dataInput_38),
    .io_dataInput_39(multiHotPriortyReductionTree_io_dataInput_39),
    .io_dataInput_40(multiHotPriortyReductionTree_io_dataInput_40),
    .io_dataInput_41(multiHotPriortyReductionTree_io_dataInput_41),
    .io_dataInput_42(multiHotPriortyReductionTree_io_dataInput_42),
    .io_dataInput_43(multiHotPriortyReductionTree_io_dataInput_43),
    .io_dataInput_44(multiHotPriortyReductionTree_io_dataInput_44),
    .io_dataInput_45(multiHotPriortyReductionTree_io_dataInput_45),
    .io_dataInput_46(multiHotPriortyReductionTree_io_dataInput_46),
    .io_dataInput_47(multiHotPriortyReductionTree_io_dataInput_47),
    .io_dataInput_48(multiHotPriortyReductionTree_io_dataInput_48),
    .io_dataInput_49(multiHotPriortyReductionTree_io_dataInput_49),
    .io_dataInput_50(multiHotPriortyReductionTree_io_dataInput_50),
    .io_dataInput_51(multiHotPriortyReductionTree_io_dataInput_51),
    .io_dataInput_52(multiHotPriortyReductionTree_io_dataInput_52),
    .io_dataInput_53(multiHotPriortyReductionTree_io_dataInput_53),
    .io_dataInput_54(multiHotPriortyReductionTree_io_dataInput_54),
    .io_dataInput_55(multiHotPriortyReductionTree_io_dataInput_55),
    .io_dataInput_56(multiHotPriortyReductionTree_io_dataInput_56),
    .io_dataInput_57(multiHotPriortyReductionTree_io_dataInput_57),
    .io_dataInput_58(multiHotPriortyReductionTree_io_dataInput_58),
    .io_dataInput_59(multiHotPriortyReductionTree_io_dataInput_59),
    .io_dataInput_60(multiHotPriortyReductionTree_io_dataInput_60),
    .io_dataInput_61(multiHotPriortyReductionTree_io_dataInput_61),
    .io_dataInput_62(multiHotPriortyReductionTree_io_dataInput_62),
    .io_dataInput_63(multiHotPriortyReductionTree_io_dataInput_63),
    .io_selectInput_0(multiHotPriortyReductionTree_io_selectInput_0),
    .io_selectInput_1(multiHotPriortyReductionTree_io_selectInput_1),
    .io_selectInput_2(multiHotPriortyReductionTree_io_selectInput_2),
    .io_selectInput_3(multiHotPriortyReductionTree_io_selectInput_3),
    .io_selectInput_4(multiHotPriortyReductionTree_io_selectInput_4),
    .io_selectInput_5(multiHotPriortyReductionTree_io_selectInput_5),
    .io_selectInput_6(multiHotPriortyReductionTree_io_selectInput_6),
    .io_selectInput_7(multiHotPriortyReductionTree_io_selectInput_7),
    .io_selectInput_8(multiHotPriortyReductionTree_io_selectInput_8),
    .io_selectInput_9(multiHotPriortyReductionTree_io_selectInput_9),
    .io_selectInput_10(multiHotPriortyReductionTree_io_selectInput_10),
    .io_selectInput_11(multiHotPriortyReductionTree_io_selectInput_11),
    .io_selectInput_12(multiHotPriortyReductionTree_io_selectInput_12),
    .io_selectInput_13(multiHotPriortyReductionTree_io_selectInput_13),
    .io_selectInput_14(multiHotPriortyReductionTree_io_selectInput_14),
    .io_selectInput_15(multiHotPriortyReductionTree_io_selectInput_15),
    .io_selectInput_16(multiHotPriortyReductionTree_io_selectInput_16),
    .io_selectInput_17(multiHotPriortyReductionTree_io_selectInput_17),
    .io_selectInput_18(multiHotPriortyReductionTree_io_selectInput_18),
    .io_selectInput_19(multiHotPriortyReductionTree_io_selectInput_19),
    .io_selectInput_20(multiHotPriortyReductionTree_io_selectInput_20),
    .io_selectInput_21(multiHotPriortyReductionTree_io_selectInput_21),
    .io_selectInput_22(multiHotPriortyReductionTree_io_selectInput_22),
    .io_selectInput_23(multiHotPriortyReductionTree_io_selectInput_23),
    .io_selectInput_24(multiHotPriortyReductionTree_io_selectInput_24),
    .io_selectInput_25(multiHotPriortyReductionTree_io_selectInput_25),
    .io_selectInput_26(multiHotPriortyReductionTree_io_selectInput_26),
    .io_selectInput_27(multiHotPriortyReductionTree_io_selectInput_27),
    .io_selectInput_28(multiHotPriortyReductionTree_io_selectInput_28),
    .io_selectInput_29(multiHotPriortyReductionTree_io_selectInput_29),
    .io_selectInput_30(multiHotPriortyReductionTree_io_selectInput_30),
    .io_selectInput_31(multiHotPriortyReductionTree_io_selectInput_31),
    .io_selectInput_32(multiHotPriortyReductionTree_io_selectInput_32),
    .io_selectInput_33(multiHotPriortyReductionTree_io_selectInput_33),
    .io_selectInput_34(multiHotPriortyReductionTree_io_selectInput_34),
    .io_selectInput_35(multiHotPriortyReductionTree_io_selectInput_35),
    .io_selectInput_36(multiHotPriortyReductionTree_io_selectInput_36),
    .io_selectInput_37(multiHotPriortyReductionTree_io_selectInput_37),
    .io_selectInput_38(multiHotPriortyReductionTree_io_selectInput_38),
    .io_selectInput_39(multiHotPriortyReductionTree_io_selectInput_39),
    .io_selectInput_40(multiHotPriortyReductionTree_io_selectInput_40),
    .io_selectInput_41(multiHotPriortyReductionTree_io_selectInput_41),
    .io_selectInput_42(multiHotPriortyReductionTree_io_selectInput_42),
    .io_selectInput_43(multiHotPriortyReductionTree_io_selectInput_43),
    .io_selectInput_44(multiHotPriortyReductionTree_io_selectInput_44),
    .io_selectInput_45(multiHotPriortyReductionTree_io_selectInput_45),
    .io_selectInput_46(multiHotPriortyReductionTree_io_selectInput_46),
    .io_selectInput_47(multiHotPriortyReductionTree_io_selectInput_47),
    .io_selectInput_48(multiHotPriortyReductionTree_io_selectInput_48),
    .io_selectInput_49(multiHotPriortyReductionTree_io_selectInput_49),
    .io_selectInput_50(multiHotPriortyReductionTree_io_selectInput_50),
    .io_selectInput_51(multiHotPriortyReductionTree_io_selectInput_51),
    .io_selectInput_52(multiHotPriortyReductionTree_io_selectInput_52),
    .io_selectInput_53(multiHotPriortyReductionTree_io_selectInput_53),
    .io_selectInput_54(multiHotPriortyReductionTree_io_selectInput_54),
    .io_selectInput_55(multiHotPriortyReductionTree_io_selectInput_55),
    .io_selectInput_56(multiHotPriortyReductionTree_io_selectInput_56),
    .io_selectInput_57(multiHotPriortyReductionTree_io_selectInput_57),
    .io_selectInput_58(multiHotPriortyReductionTree_io_selectInput_58),
    .io_selectInput_59(multiHotPriortyReductionTree_io_selectInput_59),
    .io_selectInput_60(multiHotPriortyReductionTree_io_selectInput_60),
    .io_selectInput_61(multiHotPriortyReductionTree_io_selectInput_61),
    .io_selectInput_62(multiHotPriortyReductionTree_io_selectInput_62),
    .io_selectInput_63(multiHotPriortyReductionTree_io_selectInput_63),
    .io_dataOutput(multiHotPriortyReductionTree_io_dataOutput),
    .io_selectOutput(multiHotPriortyReductionTree_io_selectOutput)
  );
  assign io_newFrame = run & _GEN_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13 71:15]
  assign io_missingFrameError = missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 131:24]
  assign io_viewBoxOutOfRangeError = viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 133:29]
  assign io_vgaRed = io_vgaRed_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 349:13]
  assign io_vgaBlue = io_vgaBlue_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 351:14]
  assign io_vgaGreen = io_vgaGreen_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 350:15]
  assign io_Hsync = io_Hsync_pipeReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 94:12]
  assign io_Vsync = io_Vsync_pipeReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 95:12]
  assign backTileMemories_0_clock = clock;
  assign backTileMemories_0_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_1_clock = clock;
  assign backTileMemories_1_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_2_clock = clock;
  assign backTileMemories_2_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_3_clock = clock;
  assign backTileMemories_3_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_4_clock = clock;
  assign backTileMemories_4_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_5_clock = clock;
  assign backTileMemories_5_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_6_clock = clock;
  assign backTileMemories_6_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_7_clock = clock;
  assign backTileMemories_7_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_8_clock = clock;
  assign backTileMemories_8_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_9_clock = clock;
  assign backTileMemories_9_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_10_clock = clock;
  assign backTileMemories_10_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_11_clock = clock;
  assign backTileMemories_11_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_12_clock = clock;
  assign backTileMemories_12_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_13_clock = clock;
  assign backTileMemories_13_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_14_clock = clock;
  assign backTileMemories_14_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_15_clock = clock;
  assign backTileMemories_15_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_16_clock = clock;
  assign backTileMemories_16_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_17_clock = clock;
  assign backTileMemories_17_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_18_clock = clock;
  assign backTileMemories_18_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_19_clock = clock;
  assign backTileMemories_19_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_20_clock = clock;
  assign backTileMemories_20_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_21_clock = clock;
  assign backTileMemories_21_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_22_clock = clock;
  assign backTileMemories_22_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_23_clock = clock;
  assign backTileMemories_23_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_24_clock = clock;
  assign backTileMemories_24_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_25_clock = clock;
  assign backTileMemories_25_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_26_clock = clock;
  assign backTileMemories_26_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_27_clock = clock;
  assign backTileMemories_27_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_28_clock = clock;
  assign backTileMemories_28_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_29_clock = clock;
  assign backTileMemories_29_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_30_clock = clock;
  assign backTileMemories_30_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_31_clock = clock;
  assign backTileMemories_31_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_32_clock = clock;
  assign backTileMemories_32_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_33_clock = clock;
  assign backTileMemories_33_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_34_clock = clock;
  assign backTileMemories_34_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_35_clock = clock;
  assign backTileMemories_35_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_36_clock = clock;
  assign backTileMemories_36_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_37_clock = clock;
  assign backTileMemories_37_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_38_clock = clock;
  assign backTileMemories_38_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_39_clock = clock;
  assign backTileMemories_39_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_40_clock = clock;
  assign backTileMemories_40_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_41_clock = clock;
  assign backTileMemories_41_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_42_clock = clock;
  assign backTileMemories_42_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_43_clock = clock;
  assign backTileMemories_43_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_44_clock = clock;
  assign backTileMemories_44_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_45_clock = clock;
  assign backTileMemories_45_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_46_clock = clock;
  assign backTileMemories_46_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_47_clock = clock;
  assign backTileMemories_47_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_48_clock = clock;
  assign backTileMemories_48_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_49_clock = clock;
  assign backTileMemories_49_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_50_clock = clock;
  assign backTileMemories_50_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_51_clock = clock;
  assign backTileMemories_51_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_52_clock = clock;
  assign backTileMemories_52_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_53_clock = clock;
  assign backTileMemories_53_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_54_clock = clock;
  assign backTileMemories_54_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_55_clock = clock;
  assign backTileMemories_55_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_56_clock = clock;
  assign backTileMemories_56_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_57_clock = clock;
  assign backTileMemories_57_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_58_clock = clock;
  assign backTileMemories_58_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_59_clock = clock;
  assign backTileMemories_59_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_60_clock = clock;
  assign backTileMemories_60_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_61_clock = clock;
  assign backTileMemories_61_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_62_clock = clock;
  assign backTileMemories_62_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_63_clock = clock;
  assign backTileMemories_63_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backBufferMemory_clock = clock;
  assign backBufferMemory_io_address = _backBufferMemory_io_address_T_5[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:31]
  assign backBufferMemory_io_writeEnable = copyEnabledReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 228:35]
  assign backBufferMemory_io_dataWrite = backBufferShadowMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 229:33]
  assign backBufferShadowMemory_clock = clock;
  assign backBufferShadowMemory_io_address = restoreEnabled ? backBufferShadowMemory_io_address_REG :
    _backBufferShadowMemory_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:43]
  assign backBufferShadowMemory_io_writeEnable = restoreEnabled & backBufferShadowMemory_io_writeEnable_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:47]
  assign backBufferShadowMemory_io_dataWrite = restoreEnabled ? backBufferRestoreMemory_io_dataRead : 6'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 224:45]
  assign backBufferRestoreMemory_clock = clock;
  assign backBufferRestoreMemory_io_address = backMemoryRestoreCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 216:65]
  assign spriteMemories_0_clock = clock;
  assign spriteMemories_0_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_1_clock = clock;
  assign spriteMemories_1_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_2_clock = clock;
  assign spriteMemories_2_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_3_clock = clock;
  assign spriteMemories_3_io_address = _spriteMemories_3_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_4_clock = clock;
  assign spriteMemories_4_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_5_clock = clock;
  assign spriteMemories_5_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_6_clock = clock;
  assign spriteMemories_6_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_7_clock = clock;
  assign spriteMemories_7_io_address = _spriteMemories_7_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_8_clock = clock;
  assign spriteMemories_8_io_address = _spriteMemories_8_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_9_clock = clock;
  assign spriteMemories_9_io_address = _spriteMemories_9_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_10_clock = clock;
  assign spriteMemories_10_io_address = _spriteMemories_10_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_11_clock = clock;
  assign spriteMemories_11_io_address = _spriteMemories_11_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_12_clock = clock;
  assign spriteMemories_12_io_address = _spriteMemories_12_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_13_clock = clock;
  assign spriteMemories_13_io_address = _spriteMemories_13_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_14_clock = clock;
  assign spriteMemories_14_io_address = _spriteMemories_14_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_15_clock = clock;
  assign spriteMemories_15_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_16_clock = clock;
  assign spriteMemories_16_io_address = _spriteMemories_16_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_17_clock = clock;
  assign spriteMemories_17_io_address = _spriteMemories_17_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_18_clock = clock;
  assign spriteMemories_18_io_address = _spriteMemories_18_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_19_clock = clock;
  assign spriteMemories_19_io_address = _spriteMemories_19_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_20_clock = clock;
  assign spriteMemories_20_io_address = _spriteMemories_20_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_21_clock = clock;
  assign spriteMemories_21_io_address = _spriteMemories_21_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_22_clock = clock;
  assign spriteMemories_22_io_address = _spriteMemories_22_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_23_clock = clock;
  assign spriteMemories_23_io_address = _spriteMemories_23_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_24_clock = clock;
  assign spriteMemories_24_io_address = _spriteMemories_24_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_25_clock = clock;
  assign spriteMemories_25_io_address = _spriteMemories_25_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_26_clock = clock;
  assign spriteMemories_26_io_address = _spriteMemories_26_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_27_clock = clock;
  assign spriteMemories_27_io_address = _spriteMemories_27_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_28_clock = clock;
  assign spriteMemories_28_io_address = _spriteMemories_28_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_29_clock = clock;
  assign spriteMemories_29_io_address = _spriteMemories_29_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_30_clock = clock;
  assign spriteMemories_30_io_address = _spriteMemories_30_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_31_clock = clock;
  assign spriteMemories_31_io_address = _spriteMemories_31_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_32_clock = clock;
  assign spriteMemories_32_io_address = _spriteMemories_32_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_33_clock = clock;
  assign spriteMemories_33_io_address = _spriteMemories_33_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_34_clock = clock;
  assign spriteMemories_34_io_address = _spriteMemories_34_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_35_clock = clock;
  assign spriteMemories_35_io_address = _spriteMemories_35_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_36_clock = clock;
  assign spriteMemories_36_io_address = _spriteMemories_36_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_37_clock = clock;
  assign spriteMemories_37_io_address = _spriteMemories_37_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_38_clock = clock;
  assign spriteMemories_38_io_address = _spriteMemories_38_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_39_clock = clock;
  assign spriteMemories_39_io_address = _spriteMemories_39_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_40_clock = clock;
  assign spriteMemories_40_io_address = _spriteMemories_40_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_41_clock = clock;
  assign spriteMemories_41_io_address = _spriteMemories_41_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_42_clock = clock;
  assign spriteMemories_42_io_address = _spriteMemories_42_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_43_clock = clock;
  assign spriteMemories_43_io_address = _spriteMemories_43_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_44_clock = clock;
  assign spriteMemories_44_io_address = _spriteMemories_44_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_45_clock = clock;
  assign spriteMemories_45_io_address = _spriteMemories_45_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_46_clock = clock;
  assign spriteMemories_46_io_address = _spriteMemories_46_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_47_clock = clock;
  assign spriteMemories_47_io_address = _spriteMemories_47_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_48_clock = clock;
  assign spriteMemories_48_io_address = _spriteMemories_48_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_49_clock = clock;
  assign spriteMemories_49_io_address = _spriteMemories_49_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_50_clock = clock;
  assign spriteMemories_50_io_address = _spriteMemories_50_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_51_clock = clock;
  assign spriteMemories_51_io_address = _spriteMemories_51_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_52_clock = clock;
  assign spriteMemories_52_io_address = _spriteMemories_52_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_53_clock = clock;
  assign spriteMemories_53_io_address = _spriteMemories_53_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_54_clock = clock;
  assign spriteMemories_54_io_address = _spriteMemories_54_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_55_clock = clock;
  assign spriteMemories_55_io_address = _spriteMemories_55_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_56_clock = clock;
  assign spriteMemories_56_io_address = _spriteMemories_56_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_57_clock = clock;
  assign spriteMemories_57_io_address = _spriteMemories_57_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_58_clock = clock;
  assign spriteMemories_58_io_address = _spriteMemories_58_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_59_clock = clock;
  assign spriteMemories_59_io_address = _spriteMemories_59_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_60_clock = clock;
  assign spriteMemories_60_io_address = _spriteMemories_60_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_61_clock = clock;
  assign spriteMemories_61_io_address = _spriteMemories_61_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_62_clock = clock;
  assign spriteMemories_62_io_address = _spriteMemories_62_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_63_clock = clock;
  assign spriteMemories_63_io_address = _spriteMemories_63_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign multiHotPriortyReductionTree_io_dataInput_0 = multiHotPriortyReductionTree_io_dataInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_1 = multiHotPriortyReductionTree_io_dataInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_2 = multiHotPriortyReductionTree_io_dataInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_3 = multiHotPriortyReductionTree_io_dataInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_4 = multiHotPriortyReductionTree_io_dataInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_5 = multiHotPriortyReductionTree_io_dataInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_6 = multiHotPriortyReductionTree_io_dataInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_7 = multiHotPriortyReductionTree_io_dataInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_8 = multiHotPriortyReductionTree_io_dataInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_9 = multiHotPriortyReductionTree_io_dataInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_10 = multiHotPriortyReductionTree_io_dataInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_11 = multiHotPriortyReductionTree_io_dataInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_12 = multiHotPriortyReductionTree_io_dataInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_13 = multiHotPriortyReductionTree_io_dataInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_14 = multiHotPriortyReductionTree_io_dataInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_15 = multiHotPriortyReductionTree_io_dataInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_16 = multiHotPriortyReductionTree_io_dataInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_17 = multiHotPriortyReductionTree_io_dataInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_18 = multiHotPriortyReductionTree_io_dataInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_19 = multiHotPriortyReductionTree_io_dataInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_20 = multiHotPriortyReductionTree_io_dataInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_21 = multiHotPriortyReductionTree_io_dataInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_22 = multiHotPriortyReductionTree_io_dataInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_23 = multiHotPriortyReductionTree_io_dataInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_24 = multiHotPriortyReductionTree_io_dataInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_25 = multiHotPriortyReductionTree_io_dataInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_26 = multiHotPriortyReductionTree_io_dataInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_27 = multiHotPriortyReductionTree_io_dataInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_28 = multiHotPriortyReductionTree_io_dataInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_29 = multiHotPriortyReductionTree_io_dataInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_30 = multiHotPriortyReductionTree_io_dataInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_31 = multiHotPriortyReductionTree_io_dataInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_32 = multiHotPriortyReductionTree_io_dataInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_33 = multiHotPriortyReductionTree_io_dataInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_34 = multiHotPriortyReductionTree_io_dataInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_35 = multiHotPriortyReductionTree_io_dataInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_36 = multiHotPriortyReductionTree_io_dataInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_37 = multiHotPriortyReductionTree_io_dataInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_38 = multiHotPriortyReductionTree_io_dataInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_39 = multiHotPriortyReductionTree_io_dataInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_40 = multiHotPriortyReductionTree_io_dataInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_41 = multiHotPriortyReductionTree_io_dataInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_42 = multiHotPriortyReductionTree_io_dataInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_43 = multiHotPriortyReductionTree_io_dataInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_44 = multiHotPriortyReductionTree_io_dataInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_45 = multiHotPriortyReductionTree_io_dataInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_46 = multiHotPriortyReductionTree_io_dataInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_47 = multiHotPriortyReductionTree_io_dataInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_48 = multiHotPriortyReductionTree_io_dataInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_49 = multiHotPriortyReductionTree_io_dataInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_50 = multiHotPriortyReductionTree_io_dataInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_51 = multiHotPriortyReductionTree_io_dataInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_52 = multiHotPriortyReductionTree_io_dataInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_53 = multiHotPriortyReductionTree_io_dataInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_54 = multiHotPriortyReductionTree_io_dataInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_55 = multiHotPriortyReductionTree_io_dataInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_56 = multiHotPriortyReductionTree_io_dataInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_57 = multiHotPriortyReductionTree_io_dataInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_58 = multiHotPriortyReductionTree_io_dataInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_59 = multiHotPriortyReductionTree_io_dataInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_60 = multiHotPriortyReductionTree_io_dataInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_61 = multiHotPriortyReductionTree_io_dataInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_62 = multiHotPriortyReductionTree_io_dataInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_63 = multiHotPriortyReductionTree_io_dataInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_selectInput_0 = multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_1 = multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_2 = multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_3 = multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_4 = multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_5 = multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_6 = multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_7 = multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_8 = multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_9 = multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_10 = multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_11 = multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_12 = multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_13 = multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_14 = multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_15 = multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_16 = multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_17 = multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_18 = multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_19 = multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_20 = multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_21 = multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_22 = multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_23 = multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_24 = multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_25 = multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_26 = multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_27 = multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_28 = multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_29 = multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_30 = multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_31 = multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_32 = multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_33 = multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_34 = multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_35 = multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_36 = multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_37 = multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_38 = multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_39 = multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_40 = multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_41 = multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_42 = multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_43 = multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_44 = multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_45 = multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_46 = multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_47 = multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_48 = multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_49 = multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_50 = multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_51 = multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_52 = multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_53 = multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_54 = multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_55 = multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_56 = multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_57 = multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_58 = multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_59 = multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_60 = multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_61 = multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_62 = multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_63 = multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
      ScaleCounterReg <= 2'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        ScaleCounterReg <= 2'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 75:23]
      end else begin
        ScaleCounterReg <= _ScaleCounterReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 88:23]
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
      CounterXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        if (CounterXReg == 10'h31f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129]
          CounterXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 77:21]
        end else begin
          CounterXReg <= _CounterXReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 85:21]
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
      CounterYReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        if (CounterXReg == 10'h31f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129]
          CounterYReg <= _GEN_0;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
      backMemoryRestoreCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
    end else if (restoreEnabled) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:70]
      backMemoryRestoreCounter <= _backMemoryRestoreCounter_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 206:30]
    end
    io_Hsync_pipeReg_0 <= io_Hsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_1 <= io_Hsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_2 <= io_Hsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_3 <= ~Hsync; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 94:27]
    io_Vsync_pipeReg_0 <= io_Vsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_1 <= io_Vsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_2 <= io_Vsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_3 <= ~Vsync; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 95:27]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
      frameClockCount <= 21'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
    end else if (frameClockCount == 21'h19a27f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 105:25]
      frameClockCount <= 21'h0;
    end else begin
      frameClockCount <= _frameClockCount_T_2;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_3 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_3 <= io_spriteXPosition_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_7 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_7 <= io_spriteXPosition_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_8 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_8 <= io_spriteXPosition_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_9 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_9 <= io_spriteXPosition_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_10 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_10 <= io_spriteXPosition_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_11 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_11 <= io_spriteXPosition_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_12 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_12 <= io_spriteXPosition_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_13 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_13 <= io_spriteXPosition_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_14 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_14 <= io_spriteXPosition_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_16 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_16 <= io_spriteXPosition_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_17 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_17 <= io_spriteXPosition_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_18 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_18 <= io_spriteXPosition_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_19 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_19 <= io_spriteXPosition_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_20 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_20 <= io_spriteXPosition_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_21 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_21 <= io_spriteXPosition_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_22 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_22 <= io_spriteXPosition_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_23 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_23 <= io_spriteXPosition_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_24 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_24 <= io_spriteXPosition_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_25 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_25 <= io_spriteXPosition_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_26 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_26 <= io_spriteXPosition_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_27 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_27 <= io_spriteXPosition_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_28 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_28 <= io_spriteXPosition_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_29 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_29 <= io_spriteXPosition_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_30 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_30 <= io_spriteXPosition_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_31 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_31 <= io_spriteXPosition_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_32 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_32 <= io_spriteXPosition_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_33 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_33 <= io_spriteXPosition_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_34 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_34 <= io_spriteXPosition_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_35 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_35 <= io_spriteXPosition_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_36 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_36 <= io_spriteXPosition_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_37 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_37 <= io_spriteXPosition_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_38 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_38 <= io_spriteXPosition_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_39 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_39 <= io_spriteXPosition_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_40 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_40 <= io_spriteXPosition_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_41 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_41 <= io_spriteXPosition_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_42 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_42 <= io_spriteXPosition_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_43 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_43 <= io_spriteXPosition_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_44 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_44 <= io_spriteXPosition_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_45 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_45 <= io_spriteXPosition_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_46 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_46 <= io_spriteXPosition_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_47 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_47 <= io_spriteXPosition_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_48 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_48 <= io_spriteXPosition_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_49 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_49 <= io_spriteXPosition_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_50 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_50 <= io_spriteXPosition_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_51 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_51 <= io_spriteXPosition_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_52 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_52 <= io_spriteXPosition_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_53 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_53 <= io_spriteXPosition_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_54 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_54 <= io_spriteXPosition_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_55 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_55 <= io_spriteXPosition_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_56 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_56 <= io_spriteXPosition_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_57 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_57 <= io_spriteXPosition_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_58 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_58 <= io_spriteXPosition_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_59 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_59 <= io_spriteXPosition_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_60 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_60 <= io_spriteXPosition_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_61 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_61 <= io_spriteXPosition_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_62 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_62 <= io_spriteXPosition_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_63 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_63 <= io_spriteXPosition_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_3 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_3 <= io_spriteYPosition_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_7 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_7 <= io_spriteYPosition_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_8 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_8 <= io_spriteYPosition_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_9 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_9 <= io_spriteYPosition_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_10 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_10 <= io_spriteYPosition_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_11 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_11 <= io_spriteYPosition_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_12 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_12 <= io_spriteYPosition_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_13 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_13 <= io_spriteYPosition_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_14 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_14 <= io_spriteYPosition_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_16 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_16 <= io_spriteYPosition_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_17 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_17 <= io_spriteYPosition_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_18 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_18 <= io_spriteYPosition_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_19 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_19 <= io_spriteYPosition_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_20 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_20 <= io_spriteYPosition_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_21 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_21 <= io_spriteYPosition_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_22 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_22 <= io_spriteYPosition_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_23 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_23 <= io_spriteYPosition_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_24 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_24 <= io_spriteYPosition_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_25 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_25 <= io_spriteYPosition_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_26 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_26 <= io_spriteYPosition_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_27 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_27 <= io_spriteYPosition_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_28 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_28 <= io_spriteYPosition_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_29 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_29 <= io_spriteYPosition_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_30 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_30 <= io_spriteYPosition_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_31 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_31 <= io_spriteYPosition_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_32 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_32 <= io_spriteYPosition_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_33 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_33 <= io_spriteYPosition_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_34 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_34 <= io_spriteYPosition_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_35 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_35 <= io_spriteYPosition_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_36 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_36 <= io_spriteYPosition_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_37 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_37 <= io_spriteYPosition_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_38 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_38 <= io_spriteYPosition_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_39 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_39 <= io_spriteYPosition_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_40 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_40 <= io_spriteYPosition_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_41 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_41 <= io_spriteYPosition_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_42 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_42 <= io_spriteYPosition_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_43 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_43 <= io_spriteYPosition_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_44 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_44 <= io_spriteYPosition_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_45 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_45 <= io_spriteYPosition_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_46 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_46 <= io_spriteYPosition_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_47 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_47 <= io_spriteYPosition_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_48 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_48 <= io_spriteYPosition_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_49 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_49 <= io_spriteYPosition_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_50 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_50 <= io_spriteYPosition_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_51 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_51 <= io_spriteYPosition_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_52 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_52 <= io_spriteYPosition_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_53 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_53 <= io_spriteYPosition_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_54 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_54 <= io_spriteYPosition_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_55 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_55 <= io_spriteYPosition_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_56 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_56 <= io_spriteYPosition_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_57 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_57 <= io_spriteYPosition_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_58 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_58 <= io_spriteYPosition_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_59 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_59 <= io_spriteYPosition_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_60 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_60 <= io_spriteYPosition_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_61 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_61 <= io_spriteYPosition_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_62 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_62 <= io_spriteYPosition_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_63 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_63 <= io_spriteYPosition_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    spriteVisibleReg_0 <= reset | _GEN_141; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_1 <= reset | _GEN_142; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_2 <= reset | _GEN_143; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_3 <= reset | _GEN_144; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_4 <= reset | _GEN_145; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_5 <= reset | _GEN_146; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_6 <= reset | _GEN_147; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_7 <= reset | _GEN_148; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_8 <= reset | _GEN_149; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_9 <= reset | _GEN_150; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_10 <= reset | _GEN_151; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_11 <= reset | _GEN_152; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_12 <= reset | _GEN_153; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_13 <= reset | _GEN_154; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_14 <= reset | _GEN_155; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_15 <= reset | _GEN_156; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_16 <= reset | _GEN_157; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_17 <= reset | _GEN_158; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_18 <= reset | _GEN_159; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_19 <= reset | _GEN_160; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_20 <= reset | _GEN_161; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_21 <= reset | _GEN_162; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_22 <= reset | _GEN_163; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_23 <= reset | _GEN_164; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_24 <= reset | _GEN_165; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_25 <= reset | _GEN_166; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_26 <= reset | _GEN_167; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_27 <= reset | _GEN_168; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_28 <= reset | _GEN_169; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_29 <= reset | _GEN_170; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_30 <= reset | _GEN_171; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_31 <= reset | _GEN_172; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_32 <= reset | _GEN_173; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_33 <= reset | _GEN_174; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_34 <= reset | _GEN_175; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_35 <= reset | _GEN_176; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_36 <= reset | _GEN_177; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_37 <= reset | _GEN_178; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_38 <= reset | _GEN_179; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_39 <= reset | _GEN_180; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_40 <= reset | _GEN_181; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_41 <= reset | _GEN_182; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_42 <= reset | _GEN_183; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_43 <= reset | _GEN_184; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_44 <= reset | _GEN_185; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_45 <= reset | _GEN_186; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_46 <= reset | _GEN_187; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_47 <= reset | _GEN_188; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_48 <= reset | _GEN_189; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_49 <= reset | _GEN_190; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_50 <= reset | _GEN_191; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_51 <= reset | _GEN_192; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_52 <= reset | _GEN_193; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_53 <= reset | _GEN_194; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_54 <= reset | _GEN_195; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_55 <= reset | _GEN_196; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_56 <= reset | _GEN_197; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_57 <= reset | _GEN_198; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_58 <= reset | _GEN_199; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_59 <= reset | _GEN_200; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_60 <= reset | _GEN_201; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_61 <= reset | _GEN_202; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_62 <= reset | _GEN_203; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_63 <= reset | _GEN_204; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_16 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_16 <= io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_17 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_17 <= io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_18 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_18 <= io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_19 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_19 <= io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_20 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_20 <= io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_21 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_21 <= io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_22 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_22 <= io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_23 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_23 <= io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_24 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_24 <= io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_25 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_25 <= io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_26 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_26 <= io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_27 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_27 <= io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_28 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_28 <= io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_29 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_29 <= io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_30 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_30 <= io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_31 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_31 <= io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_32 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_32 <= io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_33 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_33 <= io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_34 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_34 <= io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_35 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_35 <= io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_36 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_36 <= io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_37 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_37 <= io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_38 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_38 <= io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_39 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_39 <= io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_40 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_40 <= io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_41 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_41 <= io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_42 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_42 <= io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_43 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_43 <= io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_44 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_44 <= io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_45 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_45 <= io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_58 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_58 <= io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_59 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_59 <= io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_60 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_60 <= io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_16 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_16 <= io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_17 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_17 <= io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_18 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_18 <= io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_19 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_19 <= io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_20 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_20 <= io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_21 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_21 <= io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_22 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_22 <= io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_23 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_23 <= io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_24 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_24 <= io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_25 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_25 <= io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_26 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_26 <= io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_27 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_27 <= io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_28 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_28 <= io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_29 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_29 <= io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_30 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_30 <= io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_31 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_31 <= io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_32 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_32 <= io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_33 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_33 <= io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_34 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_34 <= io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_35 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_35 <= io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_36 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_36 <= io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_37 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_37 <= io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_38 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_38 <= io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_39 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_39 <= io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_40 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_40 <= io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_41 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_41 <= io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_42 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_42 <= io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_43 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_43 <= io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_44 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_44 <= io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_45 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_45 <= io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_58 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_58 <= io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_59 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_59 <= io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_60 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_60 <= io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
      viewBoxXReg <= io_viewBoxX; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
      viewBoxYReg <= 9'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
      viewBoxYReg <= io_viewBoxY; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
      missingFrameErrorReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
    end else begin
      missingFrameErrorReg <= _GEN_594;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
      viewBoxOutOfRangeErrorReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
    end else begin
      viewBoxOutOfRangeErrorReg <= _GEN_591;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
      newFrameStikyReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
    end else if (REG) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:37]
      newFrameStikyReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 152:22]
    end else begin
      newFrameStikyReg <= _GEN_592;
    end
    REG <= io_frameUpdateDone; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:16]
    backTileMemoryDataRead_0_REG <= backTileMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_1_REG <= backTileMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_2_REG <= backTileMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_3_REG <= backTileMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_4_REG <= backTileMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_5_REG <= backTileMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_6_REG <= backTileMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_7_REG <= backTileMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_8_REG <= backTileMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_9_REG <= backTileMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_10_REG <= backTileMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_11_REG <= backTileMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_12_REG <= backTileMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_13_REG <= backTileMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_14_REG <= backTileMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_15_REG <= backTileMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_16_REG <= backTileMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_17_REG <= backTileMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_18_REG <= backTileMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_19_REG <= backTileMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_20_REG <= backTileMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_21_REG <= backTileMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_22_REG <= backTileMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_23_REG <= backTileMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_24_REG <= backTileMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_25_REG <= backTileMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_26_REG <= backTileMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_27_REG <= backTileMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_28_REG <= backTileMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_29_REG <= backTileMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_30_REG <= backTileMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_31_REG <= backTileMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_32_REG <= backTileMemories_32_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_33_REG <= backTileMemories_33_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_34_REG <= backTileMemories_34_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_35_REG <= backTileMemories_35_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_36_REG <= backTileMemories_36_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_37_REG <= backTileMemories_37_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_38_REG <= backTileMemories_38_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_39_REG <= backTileMemories_39_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_40_REG <= backTileMemories_40_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_41_REG <= backTileMemories_41_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_42_REG <= backTileMemories_42_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_43_REG <= backTileMemories_43_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_44_REG <= backTileMemories_44_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_45_REG <= backTileMemories_45_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_46_REG <= backTileMemories_46_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_47_REG <= backTileMemories_47_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_48_REG <= backTileMemories_48_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_49_REG <= backTileMemories_49_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_50_REG <= backTileMemories_50_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_51_REG <= backTileMemories_51_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_52_REG <= backTileMemories_52_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_53_REG <= backTileMemories_53_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_54_REG <= backTileMemories_54_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_55_REG <= backTileMemories_55_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_56_REG <= backTileMemories_56_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_57_REG <= backTileMemories_57_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_58_REG <= backTileMemories_58_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_59_REG <= backTileMemories_59_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_60_REG <= backTileMemories_60_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_61_REG <= backTileMemories_61_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_62_REG <= backTileMemories_62_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_63_REG <= backTileMemories_63_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
      backMemoryCopyCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
    end else if (preDisplayArea) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23]
      if (backMemoryCopyCounter < 12'h800) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 187:66]
        backMemoryCopyCounter <= _backMemoryCopyCounter_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 188:29]
      end
    end else begin
      backMemoryCopyCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 197:27]
    end
    copyEnabledReg <= preDisplayArea & _T_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23 198:17]
    backBufferShadowMemory_io_address_REG <= backMemoryRestoreCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:92]
    backBufferShadowMemory_io_writeEnable_REG <= backMemoryRestoreCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:33]
    backBufferMemory_io_address_REG <= backMemoryCopyCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:83]
    fullBackgroundColor_REG <= backBufferMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:56]
    if (fullBackgroundColor[6]) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 244:25]
      pixelColorBack <= 6'h0;
    end else begin
      pixelColorBack <= fullBackgroundColor[5:0];
    end
    multiHotPriortyReductionTree_io_dataInput_0_REG <= spriteMemories_0_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1 <= spriteVisibleReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_0_REG <= spriteMemories_0_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_1_REG <= spriteMemories_1_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1 <= spriteVisibleReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_1_REG <= spriteMemories_1_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_2_REG <= spriteMemories_2_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1 <= spriteVisibleReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_2_REG <= spriteMemories_2_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_3_REG <= spriteMemories_3_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1 <= spriteVisibleReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1 <= inSpriteHorizontal_3 & inSpriteVertical_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_3_REG <= spriteMemories_3_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_4_REG <= spriteMemories_4_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1 <= spriteVisibleReg_4; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_4_REG <= spriteMemories_4_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_5_REG <= spriteMemories_5_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1 <= spriteVisibleReg_5; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_5_REG <= spriteMemories_5_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_6_REG <= spriteMemories_6_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1 <= spriteVisibleReg_6; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_6_REG <= spriteMemories_6_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_7_REG <= spriteMemories_7_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1 <= spriteVisibleReg_7; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1 <= inSpriteHorizontal_7 & inSpriteVertical_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_7_REG <= spriteMemories_7_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_8_REG <= spriteMemories_8_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1 <= spriteVisibleReg_8; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1 <= inSpriteHorizontal_8 & inSpriteVertical_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_8_REG <= spriteMemories_8_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_9_REG <= spriteMemories_9_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1 <= spriteVisibleReg_9; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1 <= inSpriteHorizontal_9 & inSpriteVertical_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_9_REG <= spriteMemories_9_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_10_REG <= spriteMemories_10_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1 <= spriteVisibleReg_10; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1 <= inSpriteHorizontal_10 & inSpriteVertical_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_10_REG <= spriteMemories_10_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_11_REG <= spriteMemories_11_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1 <= spriteVisibleReg_11; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1 <= inSpriteHorizontal_11 & inSpriteVertical_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_11_REG <= spriteMemories_11_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_12_REG <= spriteMemories_12_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1 <= spriteVisibleReg_12; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1 <= inSpriteHorizontal_12 & inSpriteVertical_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_12_REG <= spriteMemories_12_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_13_REG <= spriteMemories_13_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1 <= spriteVisibleReg_13; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1 <= inSpriteHorizontal_13 & inSpriteVertical_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_13_REG <= spriteMemories_13_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_14_REG <= spriteMemories_14_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1 <= spriteVisibleReg_14; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1 <= inSpriteHorizontal_14 & inSpriteVertical_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_14_REG <= spriteMemories_14_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_15_REG <= spriteMemories_15_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1 <= spriteVisibleReg_15; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_15_REG <= spriteMemories_15_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_16_REG <= spriteMemories_16_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1 <= spriteVisibleReg_16; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1 <= inSpriteHorizontal_16 & inSpriteVertical_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_16_REG <= spriteMemories_16_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_17_REG <= spriteMemories_17_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1 <= spriteVisibleReg_17; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1 <= inSpriteHorizontal_17 & inSpriteVertical_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_17_REG <= spriteMemories_17_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_18_REG <= spriteMemories_18_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1 <= spriteVisibleReg_18; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1 <= inSpriteHorizontal_18 & inSpriteVertical_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_18_REG <= spriteMemories_18_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_19_REG <= spriteMemories_19_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1 <= spriteVisibleReg_19; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1 <= inSpriteHorizontal_19 & inSpriteVertical_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_19_REG <= spriteMemories_19_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_20_REG <= spriteMemories_20_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1 <= spriteVisibleReg_20; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1 <= inSpriteHorizontal_20 & inSpriteVertical_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_20_REG <= spriteMemories_20_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_21_REG <= spriteMemories_21_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1 <= spriteVisibleReg_21; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1 <= inSpriteHorizontal_21 & inSpriteVertical_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_21_REG <= spriteMemories_21_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_22_REG <= spriteMemories_22_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1 <= spriteVisibleReg_22; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1 <= inSpriteHorizontal_22 & inSpriteVertical_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_22_REG <= spriteMemories_22_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_23_REG <= spriteMemories_23_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1 <= spriteVisibleReg_23; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1 <= inSpriteHorizontal_23 & inSpriteVertical_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_23_REG <= spriteMemories_23_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_24_REG <= spriteMemories_24_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1 <= spriteVisibleReg_24; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1 <= inSpriteHorizontal_24 & inSpriteVertical_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_24_REG <= spriteMemories_24_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_25_REG <= spriteMemories_25_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1 <= spriteVisibleReg_25; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1 <= inSpriteHorizontal_25 & inSpriteVertical_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_25_REG <= spriteMemories_25_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_26_REG <= spriteMemories_26_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1 <= spriteVisibleReg_26; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1 <= inSpriteHorizontal_26 & inSpriteVertical_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_26_REG <= spriteMemories_26_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_27_REG <= spriteMemories_27_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1 <= spriteVisibleReg_27; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1 <= inSpriteHorizontal_27 & inSpriteVertical_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_27_REG <= spriteMemories_27_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_28_REG <= spriteMemories_28_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1 <= spriteVisibleReg_28; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1 <= inSpriteHorizontal_28 & inSpriteVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_28_REG <= spriteMemories_28_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_29_REG <= spriteMemories_29_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1 <= spriteVisibleReg_29; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1 <= inSpriteHorizontal_29 & inSpriteVertical_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_29_REG <= spriteMemories_29_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_30_REG <= spriteMemories_30_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1 <= spriteVisibleReg_30; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1 <= inSpriteHorizontal_30 & inSpriteVertical_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_30_REG <= spriteMemories_30_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_31_REG <= spriteMemories_31_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1 <= spriteVisibleReg_31; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1 <= inSpriteHorizontal_31 & inSpriteVertical_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_31_REG <= spriteMemories_31_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_32_REG <= spriteMemories_32_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1 <= spriteVisibleReg_32; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1 <= inSpriteHorizontal_32 & inSpriteVertical_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_32_REG <= spriteMemories_32_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_33_REG <= spriteMemories_33_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1 <= spriteVisibleReg_33; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1 <= inSpriteHorizontal_33 & inSpriteVertical_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_33_REG <= spriteMemories_33_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_34_REG <= spriteMemories_34_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1 <= spriteVisibleReg_34; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1 <= inSpriteHorizontal_34 & inSpriteVertical_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_34_REG <= spriteMemories_34_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_35_REG <= spriteMemories_35_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1 <= spriteVisibleReg_35; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1 <= inSpriteHorizontal_35 & inSpriteVertical_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_35_REG <= spriteMemories_35_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_36_REG <= spriteMemories_36_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1 <= spriteVisibleReg_36; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1 <= inSpriteHorizontal_36 & inSpriteVertical_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_36_REG <= spriteMemories_36_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_37_REG <= spriteMemories_37_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1 <= spriteVisibleReg_37; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1 <= inSpriteHorizontal_37 & inSpriteVertical_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_37_REG <= spriteMemories_37_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_38_REG <= spriteMemories_38_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1 <= spriteVisibleReg_38; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1 <= inSpriteHorizontal_38 & inSpriteVertical_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_38_REG <= spriteMemories_38_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_39_REG <= spriteMemories_39_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1 <= spriteVisibleReg_39; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1 <= inSpriteHorizontal_39 & inSpriteVertical_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_39_REG <= spriteMemories_39_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_40_REG <= spriteMemories_40_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1 <= spriteVisibleReg_40; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1 <= inSpriteHorizontal_40 & inSpriteVertical_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_40_REG <= spriteMemories_40_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_41_REG <= spriteMemories_41_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1 <= spriteVisibleReg_41; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1 <= inSpriteHorizontal_41 & inSpriteVertical_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_41_REG <= spriteMemories_41_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_42_REG <= spriteMemories_42_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1 <= spriteVisibleReg_42; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1 <= inSpriteHorizontal_42 & inSpriteVertical_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_42_REG <= spriteMemories_42_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_43_REG <= spriteMemories_43_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1 <= spriteVisibleReg_43; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1 <= inSpriteHorizontal_43 & inSpriteVertical_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_43_REG <= spriteMemories_43_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_44_REG <= spriteMemories_44_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1 <= spriteVisibleReg_44; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1 <= inSpriteHorizontal_44 & inSpriteVertical_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_44_REG <= spriteMemories_44_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_45_REG <= spriteMemories_45_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1 <= spriteVisibleReg_45; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1 <= inSpriteHorizontal_45 & inSpriteVertical_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_45_REG <= spriteMemories_45_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_46_REG <= spriteMemories_46_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1 <= spriteVisibleReg_46; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1 <= inSpriteHorizontal_46 & inSpriteVertical_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_46_REG <= spriteMemories_46_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_47_REG <= spriteMemories_47_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1 <= spriteVisibleReg_47; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1 <= inSpriteHorizontal_47 & inSpriteVertical_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_47_REG <= spriteMemories_47_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_48_REG <= spriteMemories_48_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1 <= spriteVisibleReg_48; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1 <= inSpriteHorizontal_48 & inSpriteVertical_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_48_REG <= spriteMemories_48_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_49_REG <= spriteMemories_49_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1 <= spriteVisibleReg_49; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1 <= inSpriteHorizontal_49 & inSpriteVertical_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_49_REG <= spriteMemories_49_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_50_REG <= spriteMemories_50_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1 <= spriteVisibleReg_50; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1 <= inSpriteHorizontal_50 & inSpriteVertical_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_50_REG <= spriteMemories_50_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_51_REG <= spriteMemories_51_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1 <= spriteVisibleReg_51; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1 <= inSpriteHorizontal_51 & inSpriteVertical_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_51_REG <= spriteMemories_51_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_52_REG <= spriteMemories_52_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1 <= spriteVisibleReg_52; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1 <= inSpriteHorizontal_52 & inSpriteVertical_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_52_REG <= spriteMemories_52_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_53_REG <= spriteMemories_53_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1 <= spriteVisibleReg_53; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1 <= inSpriteHorizontal_53 & inSpriteVertical_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_53_REG <= spriteMemories_53_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_54_REG <= spriteMemories_54_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1 <= spriteVisibleReg_54; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1 <= inSpriteHorizontal_54 & inSpriteVertical_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_54_REG <= spriteMemories_54_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_55_REG <= spriteMemories_55_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1 <= spriteVisibleReg_55; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1 <= inSpriteHorizontal_55 & inSpriteVertical_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_55_REG <= spriteMemories_55_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_56_REG <= spriteMemories_56_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1 <= spriteVisibleReg_56; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1 <= inSpriteHorizontal_56 & inSpriteVertical_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_56_REG <= spriteMemories_56_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_57_REG <= spriteMemories_57_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1 <= spriteVisibleReg_57; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1 <= inSpriteHorizontal_57 & inSpriteVertical_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_57_REG <= spriteMemories_57_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_58_REG <= spriteMemories_58_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1 <= spriteVisibleReg_58; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1 <= inSpriteHorizontal_58 & inSpriteVertical_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_58_REG <= spriteMemories_58_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_59_REG <= spriteMemories_59_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1 <= spriteVisibleReg_59; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1 <= inSpriteHorizontal_59 & inSpriteVertical_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_59_REG <= spriteMemories_59_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_60_REG <= spriteMemories_60_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1 <= spriteVisibleReg_60; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1 <= inSpriteHorizontal_60 & inSpriteVertical_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_60_REG <= spriteMemories_60_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_61_REG <= spriteMemories_61_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1 <= spriteVisibleReg_61; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1 <= inSpriteHorizontal_61 & inSpriteVertical_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_61_REG <= spriteMemories_61_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_62_REG <= spriteMemories_62_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1 <= spriteVisibleReg_62; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1 <= inSpriteHorizontal_62 & inSpriteVertical_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_62_REG <= spriteMemories_62_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_63_REG <= spriteMemories_63_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1 <= spriteVisibleReg_63; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1 <= inSpriteHorizontal_63 & inSpriteVertical_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_63_REG <= spriteMemories_63_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    pixelColorSprite <= multiHotPriortyReductionTree_io_dataOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 339:33]
    pixelColorSpriteValid <= multiHotPriortyReductionTree_io_selectOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 340:38]
    pixelColourVGA_pipeReg_0 <= pixelColourVGA_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    pixelColourVGA_pipeReg_1 <= pixelColourVGA_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    pixelColourVGA_pipeReg_2 <= CounterXReg < 10'h280 & CounterYReg < 10'h1e0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 97:60]
    io_vgaRed_REG <= {pixelColourVGA[5:4],pixelColourVGA[5:4]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 346:26]
    io_vgaGreen_REG <= {pixelColourVGA[3:2],pixelColourVGA[3:2]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 347:28]
    io_vgaBlue_REG <= {pixelColourVGA[1:0],pixelColourVGA[1:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 348:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ScaleCounterReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  CounterXReg = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  CounterYReg = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  backMemoryRestoreCounter = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  io_Hsync_pipeReg_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_Hsync_pipeReg_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_Hsync_pipeReg_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_Hsync_pipeReg_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_Vsync_pipeReg_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  io_Vsync_pipeReg_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_Vsync_pipeReg_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_Vsync_pipeReg_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  frameClockCount = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXPositionReg_3 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXPositionReg_7 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXPositionReg_8 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXPositionReg_9 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXPositionReg_10 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXPositionReg_11 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXPositionReg_12 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteXPositionReg_13 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  spriteXPositionReg_14 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  spriteXPositionReg_16 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  spriteXPositionReg_17 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  spriteXPositionReg_18 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  spriteXPositionReg_19 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  spriteXPositionReg_20 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  spriteXPositionReg_21 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  spriteXPositionReg_22 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  spriteXPositionReg_23 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  spriteXPositionReg_24 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  spriteXPositionReg_25 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  spriteXPositionReg_26 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  spriteXPositionReg_27 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  spriteXPositionReg_28 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  spriteXPositionReg_29 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  spriteXPositionReg_30 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  spriteXPositionReg_31 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  spriteXPositionReg_32 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  spriteXPositionReg_33 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  spriteXPositionReg_34 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  spriteXPositionReg_35 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  spriteXPositionReg_36 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  spriteXPositionReg_37 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  spriteXPositionReg_38 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  spriteXPositionReg_39 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  spriteXPositionReg_40 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  spriteXPositionReg_41 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  spriteXPositionReg_42 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  spriteXPositionReg_43 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  spriteXPositionReg_44 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  spriteXPositionReg_45 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  spriteXPositionReg_46 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  spriteXPositionReg_47 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  spriteXPositionReg_48 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  spriteXPositionReg_49 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  spriteXPositionReg_50 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  spriteXPositionReg_51 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  spriteXPositionReg_52 = _RAND_58[10:0];
  _RAND_59 = {1{`RANDOM}};
  spriteXPositionReg_53 = _RAND_59[10:0];
  _RAND_60 = {1{`RANDOM}};
  spriteXPositionReg_54 = _RAND_60[10:0];
  _RAND_61 = {1{`RANDOM}};
  spriteXPositionReg_55 = _RAND_61[10:0];
  _RAND_62 = {1{`RANDOM}};
  spriteXPositionReg_56 = _RAND_62[10:0];
  _RAND_63 = {1{`RANDOM}};
  spriteXPositionReg_57 = _RAND_63[10:0];
  _RAND_64 = {1{`RANDOM}};
  spriteXPositionReg_58 = _RAND_64[10:0];
  _RAND_65 = {1{`RANDOM}};
  spriteXPositionReg_59 = _RAND_65[10:0];
  _RAND_66 = {1{`RANDOM}};
  spriteXPositionReg_60 = _RAND_66[10:0];
  _RAND_67 = {1{`RANDOM}};
  spriteXPositionReg_61 = _RAND_67[10:0];
  _RAND_68 = {1{`RANDOM}};
  spriteXPositionReg_62 = _RAND_68[10:0];
  _RAND_69 = {1{`RANDOM}};
  spriteXPositionReg_63 = _RAND_69[10:0];
  _RAND_70 = {1{`RANDOM}};
  spriteYPositionReg_3 = _RAND_70[9:0];
  _RAND_71 = {1{`RANDOM}};
  spriteYPositionReg_7 = _RAND_71[9:0];
  _RAND_72 = {1{`RANDOM}};
  spriteYPositionReg_8 = _RAND_72[9:0];
  _RAND_73 = {1{`RANDOM}};
  spriteYPositionReg_9 = _RAND_73[9:0];
  _RAND_74 = {1{`RANDOM}};
  spriteYPositionReg_10 = _RAND_74[9:0];
  _RAND_75 = {1{`RANDOM}};
  spriteYPositionReg_11 = _RAND_75[9:0];
  _RAND_76 = {1{`RANDOM}};
  spriteYPositionReg_12 = _RAND_76[9:0];
  _RAND_77 = {1{`RANDOM}};
  spriteYPositionReg_13 = _RAND_77[9:0];
  _RAND_78 = {1{`RANDOM}};
  spriteYPositionReg_14 = _RAND_78[9:0];
  _RAND_79 = {1{`RANDOM}};
  spriteYPositionReg_16 = _RAND_79[9:0];
  _RAND_80 = {1{`RANDOM}};
  spriteYPositionReg_17 = _RAND_80[9:0];
  _RAND_81 = {1{`RANDOM}};
  spriteYPositionReg_18 = _RAND_81[9:0];
  _RAND_82 = {1{`RANDOM}};
  spriteYPositionReg_19 = _RAND_82[9:0];
  _RAND_83 = {1{`RANDOM}};
  spriteYPositionReg_20 = _RAND_83[9:0];
  _RAND_84 = {1{`RANDOM}};
  spriteYPositionReg_21 = _RAND_84[9:0];
  _RAND_85 = {1{`RANDOM}};
  spriteYPositionReg_22 = _RAND_85[9:0];
  _RAND_86 = {1{`RANDOM}};
  spriteYPositionReg_23 = _RAND_86[9:0];
  _RAND_87 = {1{`RANDOM}};
  spriteYPositionReg_24 = _RAND_87[9:0];
  _RAND_88 = {1{`RANDOM}};
  spriteYPositionReg_25 = _RAND_88[9:0];
  _RAND_89 = {1{`RANDOM}};
  spriteYPositionReg_26 = _RAND_89[9:0];
  _RAND_90 = {1{`RANDOM}};
  spriteYPositionReg_27 = _RAND_90[9:0];
  _RAND_91 = {1{`RANDOM}};
  spriteYPositionReg_28 = _RAND_91[9:0];
  _RAND_92 = {1{`RANDOM}};
  spriteYPositionReg_29 = _RAND_92[9:0];
  _RAND_93 = {1{`RANDOM}};
  spriteYPositionReg_30 = _RAND_93[9:0];
  _RAND_94 = {1{`RANDOM}};
  spriteYPositionReg_31 = _RAND_94[9:0];
  _RAND_95 = {1{`RANDOM}};
  spriteYPositionReg_32 = _RAND_95[9:0];
  _RAND_96 = {1{`RANDOM}};
  spriteYPositionReg_33 = _RAND_96[9:0];
  _RAND_97 = {1{`RANDOM}};
  spriteYPositionReg_34 = _RAND_97[9:0];
  _RAND_98 = {1{`RANDOM}};
  spriteYPositionReg_35 = _RAND_98[9:0];
  _RAND_99 = {1{`RANDOM}};
  spriteYPositionReg_36 = _RAND_99[9:0];
  _RAND_100 = {1{`RANDOM}};
  spriteYPositionReg_37 = _RAND_100[9:0];
  _RAND_101 = {1{`RANDOM}};
  spriteYPositionReg_38 = _RAND_101[9:0];
  _RAND_102 = {1{`RANDOM}};
  spriteYPositionReg_39 = _RAND_102[9:0];
  _RAND_103 = {1{`RANDOM}};
  spriteYPositionReg_40 = _RAND_103[9:0];
  _RAND_104 = {1{`RANDOM}};
  spriteYPositionReg_41 = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  spriteYPositionReg_42 = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  spriteYPositionReg_43 = _RAND_106[9:0];
  _RAND_107 = {1{`RANDOM}};
  spriteYPositionReg_44 = _RAND_107[9:0];
  _RAND_108 = {1{`RANDOM}};
  spriteYPositionReg_45 = _RAND_108[9:0];
  _RAND_109 = {1{`RANDOM}};
  spriteYPositionReg_46 = _RAND_109[9:0];
  _RAND_110 = {1{`RANDOM}};
  spriteYPositionReg_47 = _RAND_110[9:0];
  _RAND_111 = {1{`RANDOM}};
  spriteYPositionReg_48 = _RAND_111[9:0];
  _RAND_112 = {1{`RANDOM}};
  spriteYPositionReg_49 = _RAND_112[9:0];
  _RAND_113 = {1{`RANDOM}};
  spriteYPositionReg_50 = _RAND_113[9:0];
  _RAND_114 = {1{`RANDOM}};
  spriteYPositionReg_51 = _RAND_114[9:0];
  _RAND_115 = {1{`RANDOM}};
  spriteYPositionReg_52 = _RAND_115[9:0];
  _RAND_116 = {1{`RANDOM}};
  spriteYPositionReg_53 = _RAND_116[9:0];
  _RAND_117 = {1{`RANDOM}};
  spriteYPositionReg_54 = _RAND_117[9:0];
  _RAND_118 = {1{`RANDOM}};
  spriteYPositionReg_55 = _RAND_118[9:0];
  _RAND_119 = {1{`RANDOM}};
  spriteYPositionReg_56 = _RAND_119[9:0];
  _RAND_120 = {1{`RANDOM}};
  spriteYPositionReg_57 = _RAND_120[9:0];
  _RAND_121 = {1{`RANDOM}};
  spriteYPositionReg_58 = _RAND_121[9:0];
  _RAND_122 = {1{`RANDOM}};
  spriteYPositionReg_59 = _RAND_122[9:0];
  _RAND_123 = {1{`RANDOM}};
  spriteYPositionReg_60 = _RAND_123[9:0];
  _RAND_124 = {1{`RANDOM}};
  spriteYPositionReg_61 = _RAND_124[9:0];
  _RAND_125 = {1{`RANDOM}};
  spriteYPositionReg_62 = _RAND_125[9:0];
  _RAND_126 = {1{`RANDOM}};
  spriteYPositionReg_63 = _RAND_126[9:0];
  _RAND_127 = {1{`RANDOM}};
  spriteVisibleReg_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  spriteVisibleReg_1 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  spriteVisibleReg_2 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  spriteVisibleReg_3 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  spriteVisibleReg_4 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  spriteVisibleReg_5 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  spriteVisibleReg_6 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  spriteVisibleReg_7 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  spriteVisibleReg_8 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  spriteVisibleReg_9 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  spriteVisibleReg_10 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  spriteVisibleReg_11 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  spriteVisibleReg_12 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  spriteVisibleReg_13 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  spriteVisibleReg_14 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  spriteVisibleReg_15 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  spriteVisibleReg_16 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  spriteVisibleReg_17 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  spriteVisibleReg_18 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  spriteVisibleReg_19 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  spriteVisibleReg_20 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  spriteVisibleReg_21 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  spriteVisibleReg_22 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  spriteVisibleReg_23 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  spriteVisibleReg_24 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  spriteVisibleReg_25 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  spriteVisibleReg_26 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  spriteVisibleReg_27 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  spriteVisibleReg_28 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  spriteVisibleReg_29 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  spriteVisibleReg_30 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  spriteVisibleReg_31 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  spriteVisibleReg_32 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  spriteVisibleReg_33 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  spriteVisibleReg_34 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  spriteVisibleReg_35 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  spriteVisibleReg_36 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  spriteVisibleReg_37 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  spriteVisibleReg_38 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  spriteVisibleReg_39 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  spriteVisibleReg_40 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  spriteVisibleReg_41 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  spriteVisibleReg_42 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  spriteVisibleReg_43 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  spriteVisibleReg_44 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  spriteVisibleReg_45 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  spriteVisibleReg_46 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  spriteVisibleReg_47 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  spriteVisibleReg_48 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  spriteVisibleReg_49 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  spriteVisibleReg_50 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  spriteVisibleReg_51 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  spriteVisibleReg_52 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  spriteVisibleReg_53 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  spriteVisibleReg_54 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  spriteVisibleReg_55 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  spriteVisibleReg_56 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  spriteVisibleReg_57 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  spriteVisibleReg_58 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  spriteVisibleReg_59 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  spriteVisibleReg_60 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  spriteVisibleReg_61 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  spriteVisibleReg_62 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  spriteVisibleReg_63 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_16 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_17 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_18 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_19 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_20 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_21 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_22 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_23 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_24 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_25 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_26 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_27 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_28 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_29 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_30 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_31 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_32 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_33 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_34 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_35 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_36 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_37 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_38 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_39 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_40 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_41 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_42 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_43 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_44 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_45 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_58 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_59 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_60 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_16 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_17 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_18 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_19 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_20 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_21 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_22 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_23 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_24 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_25 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_26 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_27 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_28 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_29 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_30 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_31 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_32 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_33 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_34 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_35 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_36 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_37 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_38 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_39 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_40 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_41 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_42 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_43 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_44 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_45 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_58 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_59 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_60 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  viewBoxXReg = _RAND_257[9:0];
  _RAND_258 = {1{`RANDOM}};
  viewBoxYReg = _RAND_258[8:0];
  _RAND_259 = {1{`RANDOM}};
  missingFrameErrorReg = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  viewBoxOutOfRangeErrorReg = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  newFrameStikyReg = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  REG = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  backTileMemoryDataRead_0_REG = _RAND_263[6:0];
  _RAND_264 = {1{`RANDOM}};
  backTileMemoryDataRead_1_REG = _RAND_264[6:0];
  _RAND_265 = {1{`RANDOM}};
  backTileMemoryDataRead_2_REG = _RAND_265[6:0];
  _RAND_266 = {1{`RANDOM}};
  backTileMemoryDataRead_3_REG = _RAND_266[6:0];
  _RAND_267 = {1{`RANDOM}};
  backTileMemoryDataRead_4_REG = _RAND_267[6:0];
  _RAND_268 = {1{`RANDOM}};
  backTileMemoryDataRead_5_REG = _RAND_268[6:0];
  _RAND_269 = {1{`RANDOM}};
  backTileMemoryDataRead_6_REG = _RAND_269[6:0];
  _RAND_270 = {1{`RANDOM}};
  backTileMemoryDataRead_7_REG = _RAND_270[6:0];
  _RAND_271 = {1{`RANDOM}};
  backTileMemoryDataRead_8_REG = _RAND_271[6:0];
  _RAND_272 = {1{`RANDOM}};
  backTileMemoryDataRead_9_REG = _RAND_272[6:0];
  _RAND_273 = {1{`RANDOM}};
  backTileMemoryDataRead_10_REG = _RAND_273[6:0];
  _RAND_274 = {1{`RANDOM}};
  backTileMemoryDataRead_11_REG = _RAND_274[6:0];
  _RAND_275 = {1{`RANDOM}};
  backTileMemoryDataRead_12_REG = _RAND_275[6:0];
  _RAND_276 = {1{`RANDOM}};
  backTileMemoryDataRead_13_REG = _RAND_276[6:0];
  _RAND_277 = {1{`RANDOM}};
  backTileMemoryDataRead_14_REG = _RAND_277[6:0];
  _RAND_278 = {1{`RANDOM}};
  backTileMemoryDataRead_15_REG = _RAND_278[6:0];
  _RAND_279 = {1{`RANDOM}};
  backTileMemoryDataRead_16_REG = _RAND_279[6:0];
  _RAND_280 = {1{`RANDOM}};
  backTileMemoryDataRead_17_REG = _RAND_280[6:0];
  _RAND_281 = {1{`RANDOM}};
  backTileMemoryDataRead_18_REG = _RAND_281[6:0];
  _RAND_282 = {1{`RANDOM}};
  backTileMemoryDataRead_19_REG = _RAND_282[6:0];
  _RAND_283 = {1{`RANDOM}};
  backTileMemoryDataRead_20_REG = _RAND_283[6:0];
  _RAND_284 = {1{`RANDOM}};
  backTileMemoryDataRead_21_REG = _RAND_284[6:0];
  _RAND_285 = {1{`RANDOM}};
  backTileMemoryDataRead_22_REG = _RAND_285[6:0];
  _RAND_286 = {1{`RANDOM}};
  backTileMemoryDataRead_23_REG = _RAND_286[6:0];
  _RAND_287 = {1{`RANDOM}};
  backTileMemoryDataRead_24_REG = _RAND_287[6:0];
  _RAND_288 = {1{`RANDOM}};
  backTileMemoryDataRead_25_REG = _RAND_288[6:0];
  _RAND_289 = {1{`RANDOM}};
  backTileMemoryDataRead_26_REG = _RAND_289[6:0];
  _RAND_290 = {1{`RANDOM}};
  backTileMemoryDataRead_27_REG = _RAND_290[6:0];
  _RAND_291 = {1{`RANDOM}};
  backTileMemoryDataRead_28_REG = _RAND_291[6:0];
  _RAND_292 = {1{`RANDOM}};
  backTileMemoryDataRead_29_REG = _RAND_292[6:0];
  _RAND_293 = {1{`RANDOM}};
  backTileMemoryDataRead_30_REG = _RAND_293[6:0];
  _RAND_294 = {1{`RANDOM}};
  backTileMemoryDataRead_31_REG = _RAND_294[6:0];
  _RAND_295 = {1{`RANDOM}};
  backTileMemoryDataRead_32_REG = _RAND_295[6:0];
  _RAND_296 = {1{`RANDOM}};
  backTileMemoryDataRead_33_REG = _RAND_296[6:0];
  _RAND_297 = {1{`RANDOM}};
  backTileMemoryDataRead_34_REG = _RAND_297[6:0];
  _RAND_298 = {1{`RANDOM}};
  backTileMemoryDataRead_35_REG = _RAND_298[6:0];
  _RAND_299 = {1{`RANDOM}};
  backTileMemoryDataRead_36_REG = _RAND_299[6:0];
  _RAND_300 = {1{`RANDOM}};
  backTileMemoryDataRead_37_REG = _RAND_300[6:0];
  _RAND_301 = {1{`RANDOM}};
  backTileMemoryDataRead_38_REG = _RAND_301[6:0];
  _RAND_302 = {1{`RANDOM}};
  backTileMemoryDataRead_39_REG = _RAND_302[6:0];
  _RAND_303 = {1{`RANDOM}};
  backTileMemoryDataRead_40_REG = _RAND_303[6:0];
  _RAND_304 = {1{`RANDOM}};
  backTileMemoryDataRead_41_REG = _RAND_304[6:0];
  _RAND_305 = {1{`RANDOM}};
  backTileMemoryDataRead_42_REG = _RAND_305[6:0];
  _RAND_306 = {1{`RANDOM}};
  backTileMemoryDataRead_43_REG = _RAND_306[6:0];
  _RAND_307 = {1{`RANDOM}};
  backTileMemoryDataRead_44_REG = _RAND_307[6:0];
  _RAND_308 = {1{`RANDOM}};
  backTileMemoryDataRead_45_REG = _RAND_308[6:0];
  _RAND_309 = {1{`RANDOM}};
  backTileMemoryDataRead_46_REG = _RAND_309[6:0];
  _RAND_310 = {1{`RANDOM}};
  backTileMemoryDataRead_47_REG = _RAND_310[6:0];
  _RAND_311 = {1{`RANDOM}};
  backTileMemoryDataRead_48_REG = _RAND_311[6:0];
  _RAND_312 = {1{`RANDOM}};
  backTileMemoryDataRead_49_REG = _RAND_312[6:0];
  _RAND_313 = {1{`RANDOM}};
  backTileMemoryDataRead_50_REG = _RAND_313[6:0];
  _RAND_314 = {1{`RANDOM}};
  backTileMemoryDataRead_51_REG = _RAND_314[6:0];
  _RAND_315 = {1{`RANDOM}};
  backTileMemoryDataRead_52_REG = _RAND_315[6:0];
  _RAND_316 = {1{`RANDOM}};
  backTileMemoryDataRead_53_REG = _RAND_316[6:0];
  _RAND_317 = {1{`RANDOM}};
  backTileMemoryDataRead_54_REG = _RAND_317[6:0];
  _RAND_318 = {1{`RANDOM}};
  backTileMemoryDataRead_55_REG = _RAND_318[6:0];
  _RAND_319 = {1{`RANDOM}};
  backTileMemoryDataRead_56_REG = _RAND_319[6:0];
  _RAND_320 = {1{`RANDOM}};
  backTileMemoryDataRead_57_REG = _RAND_320[6:0];
  _RAND_321 = {1{`RANDOM}};
  backTileMemoryDataRead_58_REG = _RAND_321[6:0];
  _RAND_322 = {1{`RANDOM}};
  backTileMemoryDataRead_59_REG = _RAND_322[6:0];
  _RAND_323 = {1{`RANDOM}};
  backTileMemoryDataRead_60_REG = _RAND_323[6:0];
  _RAND_324 = {1{`RANDOM}};
  backTileMemoryDataRead_61_REG = _RAND_324[6:0];
  _RAND_325 = {1{`RANDOM}};
  backTileMemoryDataRead_62_REG = _RAND_325[6:0];
  _RAND_326 = {1{`RANDOM}};
  backTileMemoryDataRead_63_REG = _RAND_326[6:0];
  _RAND_327 = {1{`RANDOM}};
  backMemoryCopyCounter = _RAND_327[11:0];
  _RAND_328 = {1{`RANDOM}};
  copyEnabledReg = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  backBufferShadowMemory_io_address_REG = _RAND_329[10:0];
  _RAND_330 = {1{`RANDOM}};
  backBufferShadowMemory_io_writeEnable_REG = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  backBufferMemory_io_address_REG = _RAND_331[10:0];
  _RAND_332 = {1{`RANDOM}};
  fullBackgroundColor_REG = _RAND_332[5:0];
  _RAND_333 = {1{`RANDOM}};
  pixelColorBack = _RAND_333[5:0];
  _RAND_334 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_0_REG = _RAND_334[5:0];
  _RAND_335 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_REG = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_1_REG = _RAND_340[5:0];
  _RAND_341 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_REG = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_2_REG = _RAND_346[5:0];
  _RAND_347 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_REG = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_3_REG = _RAND_352[5:0];
  _RAND_353 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_REG = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_4_REG = _RAND_358[5:0];
  _RAND_359 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_REG = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_5_REG = _RAND_364[5:0];
  _RAND_365 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_REG = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_6_REG = _RAND_370[5:0];
  _RAND_371 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_REG = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_7_REG = _RAND_376[5:0];
  _RAND_377 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_REG = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_8_REG = _RAND_382[5:0];
  _RAND_383 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_REG = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_9_REG = _RAND_388[5:0];
  _RAND_389 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_REG = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_10_REG = _RAND_394[5:0];
  _RAND_395 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_REG = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_11_REG = _RAND_400[5:0];
  _RAND_401 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_REG = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_12_REG = _RAND_406[5:0];
  _RAND_407 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_REG = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_13_REG = _RAND_412[5:0];
  _RAND_413 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_REG = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_14_REG = _RAND_418[5:0];
  _RAND_419 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_REG = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_15_REG = _RAND_424[5:0];
  _RAND_425 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_REG = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_16_REG = _RAND_430[5:0];
  _RAND_431 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_REG = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_17_REG = _RAND_436[5:0];
  _RAND_437 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_REG = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_18_REG = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_REG = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_19_REG = _RAND_448[5:0];
  _RAND_449 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_REG = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_20_REG = _RAND_454[5:0];
  _RAND_455 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_REG = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_21_REG = _RAND_460[5:0];
  _RAND_461 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_REG = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_22_REG = _RAND_466[5:0];
  _RAND_467 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_REG = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_23_REG = _RAND_472[5:0];
  _RAND_473 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_REG = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_24_REG = _RAND_478[5:0];
  _RAND_479 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_REG = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_25_REG = _RAND_484[5:0];
  _RAND_485 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_REG = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_26_REG = _RAND_490[5:0];
  _RAND_491 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_REG = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_27_REG = _RAND_496[5:0];
  _RAND_497 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_REG = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_28_REG = _RAND_502[5:0];
  _RAND_503 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_REG = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_29_REG = _RAND_508[5:0];
  _RAND_509 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_REG = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_30_REG = _RAND_514[5:0];
  _RAND_515 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_REG = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_31_REG = _RAND_520[5:0];
  _RAND_521 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_REG = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_32_REG = _RAND_526[5:0];
  _RAND_527 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_REG = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_33_REG = _RAND_532[5:0];
  _RAND_533 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_REG = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_34_REG = _RAND_538[5:0];
  _RAND_539 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_REG = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_35_REG = _RAND_544[5:0];
  _RAND_545 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_REG = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_36_REG = _RAND_550[5:0];
  _RAND_551 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_REG = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_37_REG = _RAND_556[5:0];
  _RAND_557 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_REG = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_38_REG = _RAND_562[5:0];
  _RAND_563 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_REG = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_39_REG = _RAND_568[5:0];
  _RAND_569 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_REG = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_40_REG = _RAND_574[5:0];
  _RAND_575 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_REG = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_41_REG = _RAND_580[5:0];
  _RAND_581 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_REG = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_42_REG = _RAND_586[5:0];
  _RAND_587 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_REG = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_43_REG = _RAND_592[5:0];
  _RAND_593 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_REG = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_44_REG = _RAND_598[5:0];
  _RAND_599 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_REG = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_45_REG = _RAND_604[5:0];
  _RAND_605 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_REG = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_46_REG = _RAND_610[5:0];
  _RAND_611 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_REG = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_47_REG = _RAND_616[5:0];
  _RAND_617 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_REG = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_48_REG = _RAND_622[5:0];
  _RAND_623 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_REG = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_49_REG = _RAND_628[5:0];
  _RAND_629 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_REG = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_50_REG = _RAND_634[5:0];
  _RAND_635 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_REG = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_51_REG = _RAND_640[5:0];
  _RAND_641 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_REG = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_52_REG = _RAND_646[5:0];
  _RAND_647 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_REG = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_53_REG = _RAND_652[5:0];
  _RAND_653 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_REG = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_54_REG = _RAND_658[5:0];
  _RAND_659 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_REG = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_55_REG = _RAND_664[5:0];
  _RAND_665 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_REG = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_56_REG = _RAND_670[5:0];
  _RAND_671 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_REG = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_57_REG = _RAND_676[5:0];
  _RAND_677 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_REG = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_58_REG = _RAND_682[5:0];
  _RAND_683 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_REG = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_59_REG = _RAND_688[5:0];
  _RAND_689 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_REG = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_60_REG = _RAND_694[5:0];
  _RAND_695 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_REG = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_61_REG = _RAND_700[5:0];
  _RAND_701 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_REG = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_62_REG = _RAND_706[5:0];
  _RAND_707 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_REG = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_63_REG = _RAND_712[5:0];
  _RAND_713 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_REG = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  pixelColorSprite = _RAND_718[5:0];
  _RAND_719 = {1{`RANDOM}};
  pixelColorSpriteValid = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_0 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_1 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_2 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  io_vgaRed_REG = _RAND_723[3:0];
  _RAND_724 = {1{`RANDOM}};
  io_vgaGreen_REG = _RAND_724[3:0];
  _RAND_725 = {1{`RANDOM}};
  io_vgaBlue_REG = _RAND_725[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Memory_131(
  input         clock,
  input  [7:0]  io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [27:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [7:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(8), .DATA_WIDTH(28), .LOAD_FILE("memory_init/tune_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 28'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_132(
  input         clock,
  input  [7:0]  io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [27:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [7:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(8), .DATA_WIDTH(28), .LOAD_FILE("memory_init/tune_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 28'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module SoundEngine(
  input   clock,
  input   reset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  tuneMemories_0_clock; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [7:0] tuneMemories_0_io_address; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [27:0] tuneMemories_0_io_dataRead; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire  tuneMemories_1_clock; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [7:0] tuneMemories_1_io_address; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [27:0] tuneMemories_1_io_dataRead; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  reg [11:0] durationCountReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
  reg [11:0] durationCountReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
  reg [11:0] currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
  reg [11:0] currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
  reg [7:0] nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
  reg [7:0] nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
  reg [1:0] stateReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
  reg [1:0] stateReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
  reg  newNoteLoadReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
  reg  newNoteLoadReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
  wire  durationCountRegDone_0 = durationCountReg_0 == 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 89:54]
  wire  _T_8 = tuneMemories_0_io_dataRead[27:16] != 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 111:60]
  wire [1:0] _GEN_4 = tuneMemories_0_io_dataRead[27:16] != 12'h0 ? 2'h3 : stateReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 112:23 62:25]
  wire [11:0] _GEN_6 = tuneMemories_0_io_dataRead[27:16] != 12'h0 ? tuneMemories_0_io_dataRead[27:16] :
    currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 114:30 58:32]
  wire  _T_13 = durationCountRegDone_0 & ~newNoteLoadReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:44]
  wire [7:0] _nextIndexReg_0_T_1 = nextIndexReg_0 + 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 126:46]
  wire [11:0] _GEN_10 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? tuneMemories_0_io_dataRead[27:16] :
    currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 124:30 58:32]
  wire [7:0] _GEN_12 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? _nextIndexReg_0_T_1 : nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 126:27 59:29]
  wire [7:0] _GEN_14 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? 8'h0 : _GEN_12; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 120:27]
  wire [11:0] _GEN_16 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? currDurationReg_0 : _GEN_10; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 58:32]
  wire  _GEN_17 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? 1'h0 : _T_13; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 97:23]
  wire [7:0] _GEN_22 = 2'h3 == stateReg_0 ? _GEN_14 : nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 59:29]
  wire [11:0] _GEN_24 = 2'h3 == stateReg_0 ? _GEN_16 : currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 58:32]
  wire  _GEN_25 = 2'h3 == stateReg_0 & _GEN_17; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 97:23]
  wire  durationCountRegDone_1 = durationCountReg_1 == 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 89:54]
  wire  _T_25 = tuneMemories_1_io_dataRead[27:16] != 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 111:60]
  wire [1:0] _GEN_52 = tuneMemories_1_io_dataRead[27:16] != 12'h0 ? 2'h3 : stateReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 112:23 62:25]
  wire [11:0] _GEN_54 = tuneMemories_1_io_dataRead[27:16] != 12'h0 ? tuneMemories_1_io_dataRead[27:16] :
    currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 114:30 58:32]
  wire  _T_30 = durationCountRegDone_1 & ~newNoteLoadReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:44]
  wire [7:0] _nextIndexReg_1_T_1 = nextIndexReg_1 + 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 126:46]
  wire [11:0] _GEN_58 = durationCountRegDone_1 & ~newNoteLoadReg_1 ? tuneMemories_1_io_dataRead[27:16] :
    currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 124:30 58:32]
  wire [7:0] _GEN_60 = durationCountRegDone_1 & ~newNoteLoadReg_1 ? _nextIndexReg_1_T_1 : nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 126:27 59:29]
  wire [7:0] _GEN_62 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? 8'h0 : _GEN_60; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 120:27]
  wire [11:0] _GEN_64 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? currDurationReg_1 : _GEN_58; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 58:32]
  wire  _GEN_65 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? 1'h0 : _T_30; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 97:23]
  wire [7:0] _GEN_70 = 2'h3 == stateReg_1 ? _GEN_62 : nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 59:29]
  wire [11:0] _GEN_72 = 2'h3 == stateReg_1 ? _GEN_64 : currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 58:32]
  wire  _GEN_73 = 2'h3 == stateReg_1 & _GEN_65; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 97:23]
  Memory_131 tuneMemories_0 ( // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
    .clock(tuneMemories_0_clock),
    .io_address(tuneMemories_0_io_address),
    .io_dataRead(tuneMemories_0_io_dataRead)
  );
  Memory_132 tuneMemories_1 ( // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
    .clock(tuneMemories_1_clock),
    .io_address(tuneMemories_1_io_address),
    .io_dataRead(tuneMemories_1_io_dataRead)
  );
  assign tuneMemories_0_clock = clock;
  assign tuneMemories_0_io_address = nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 72:32]
  assign tuneMemories_1_clock = clock;
  assign tuneMemories_1_io_address = nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 72:32]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
      durationCountReg_0 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
    end else if (newNoteLoadReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 84:35]
      durationCountReg_0 <= currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 85:27]
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
      durationCountReg_1 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
    end else if (newNoteLoadReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 84:35]
      durationCountReg_1 <= currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 85:27]
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
      currDurationReg_0 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
    end else if (!(2'h0 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h1 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
          currDurationReg_0 <= _GEN_6;
        end else begin
          currDurationReg_0 <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
      currDurationReg_1 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
    end else if (!(2'h0 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h1 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
          currDurationReg_1 <= _GEN_54;
        end else begin
          currDurationReg_1 <= _GEN_72;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
      nextIndexReg_0 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 102:25]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 107:25]
    end else if (!(2'h2 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= _GEN_22;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
      nextIndexReg_1 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 102:25]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 107:25]
    end else if (!(2'h2 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= _GEN_70;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
      stateReg_0 <= 2'h0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= 2'h1; // @[\\src\\main\\scala\\SoundEngine.scala 103:21]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= 2'h2; // @[\\src\\main\\scala\\SoundEngine.scala 108:21]
    end else if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= _GEN_4;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
      stateReg_1 <= 2'h0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= 2'h1; // @[\\src\\main\\scala\\SoundEngine.scala 103:21]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= 2'h2; // @[\\src\\main\\scala\\SoundEngine.scala 108:21]
    end else if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= _GEN_52;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= _T_8;
    end else begin
      newNoteLoadReg_0 <= _GEN_25;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= _T_25;
    end else begin
      newNoteLoadReg_1 <= _GEN_73;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  durationCountReg_0 = _RAND_0[11:0];
  _RAND_1 = {1{`RANDOM}};
  durationCountReg_1 = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  currDurationReg_0 = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  currDurationReg_1 = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  nextIndexReg_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  nextIndexReg_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  stateReg_0 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  stateReg_1 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  newNoteLoadReg_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  newNoteLoadReg_1 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Difficulty(
  input         clock,
  input         reset,
  input  [1:0]  io_level, // @[\\src\\main\\scala\\Difficulty.scala 5:14]
  output [26:0] io_speed, // @[\\src\\main\\scala\\Difficulty.scala 5:14]
  input         io_resetSpeed // @[\\src\\main\\scala\\Difficulty.scala 5:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [26:0] speedCnt; // @[\\src\\main\\scala\\Difficulty.scala 13:25]
  reg [26:0] frameDivider; // @[\\src\\main\\scala\\Difficulty.scala 16:29]
  wire  tick = frameDivider == 27'h196e6a; // @[\\src\\main\\scala\\Difficulty.scala 23:21]
  wire [26:0] _frameDivider_T_1 = frameDivider + 27'h1; // @[\\src\\main\\scala\\Difficulty.scala 27:34]
  wire [26:0] _speedCnt_T_1 = speedCnt + 27'h1; // @[\\src\\main\\scala\\Difficulty.scala 34:26]
  wire [21:0] timeInSeconds = speedCnt[26:5]; // @[\\src\\main\\scala\\Difficulty.scala 39:32]
  wire [1:0] _speedFactor_T_1 = 2'h1 == io_level ? $signed(2'sh1) : $signed(2'sh0); // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire  _speedFactor_T_2 = 2'h2 == io_level; // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [1:0] _speedFactor_T_3 = 2'h2 == io_level ? $signed(2'sh1) : $signed(_speedFactor_T_1); // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire  _speedFactor_T_4 = 2'h3 == io_level; // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [2:0] speedFactor = 2'h3 == io_level ? $signed(3'sh2) : $signed({{1{_speedFactor_T_3[1]}},_speedFactor_T_3}); // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [17:0] _rawSpeed_T = timeInSeconds[21:4]; // @[\\src\\main\\scala\\Difficulty.scala 47:36]
  wire [20:0] _rawSpeed_T_1 = $signed(_rawSpeed_T) * $signed(speedFactor); // @[\\src\\main\\scala\\Difficulty.scala 47:43]
  wire [20:0] rawSpeed = 21'sh1 + $signed(_rawSpeed_T_1); // @[\\src\\main\\scala\\Difficulty.scala 47:22]
  wire [4:0] _speedCap_T_3 = _speedFactor_T_2 ? $signed(5'shf) : $signed(5'sha); // @[\\src\\main\\scala\\Difficulty.scala 49:43]
  wire [5:0] speedCap = _speedFactor_T_4 ? $signed(6'sh14) : $signed({{1{_speedCap_T_3[4]}},_speedCap_T_3}); // @[\\src\\main\\scala\\Difficulty.scala 49:43]
  wire [20:0] _GEN_4 = {{15{speedCap[5]}},speedCap}; // @[\\src\\main\\scala\\Difficulty.scala 54:28]
  wire [20:0] _io_speed_T_1 = $signed(rawSpeed) > $signed(_GEN_4) ? $signed({{15{speedCap[5]}},speedCap}) : $signed(
    rawSpeed); // @[\\src\\main\\scala\\Difficulty.scala 54:18]
  assign io_speed = {{6{_io_speed_T_1[20]}},_io_speed_T_1}; // @[\\src\\main\\scala\\Difficulty.scala 54:12]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\Difficulty.scala 13:25]
      speedCnt <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 13:25]
    end else if (io_resetSpeed) begin // @[\\src\\main\\scala\\Difficulty.scala 31:23]
      speedCnt <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 32:14]
    end else if (tick) begin // @[\\src\\main\\scala\\Difficulty.scala 33:20]
      speedCnt <= _speedCnt_T_1; // @[\\src\\main\\scala\\Difficulty.scala 34:14]
    end
    if (reset) begin // @[\\src\\main\\scala\\Difficulty.scala 16:29]
      frameDivider <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 16:29]
    end else if (tick) begin // @[\\src\\main\\scala\\Difficulty.scala 23:37]
      frameDivider <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 24:18]
    end else begin
      frameDivider <= _frameDivider_T_1; // @[\\src\\main\\scala\\Difficulty.scala 27:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  speedCnt = _RAND_0[26:0];
  _RAND_1 = {1{`RANDOM}};
  frameDivider = _RAND_1[26:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LFSR(
  input        clock,
  input        reset,
  output [9:0] io_out_0, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_1, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_2, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_3, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_4, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_5, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_6, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_7, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_8, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_9, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_20, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_21, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_22, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_23, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_24, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_25, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_26, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_27, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_28, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_29 // @[\\src\\main\\scala\\LFSR.scala 5:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] reg_; // @[\\src\\main\\scala\\LFSR.scala 10:20]
  wire  feedback = reg_[63] ^ reg_[62] ^ reg_[60] ^ reg_[59]; // @[\\src\\main\\scala\\LFSR.scala 13:46]
  wire [63:0] _reg_T_1 = {reg_[62:0],feedback}; // @[\\src\\main\\scala\\LFSR.scala 16:13]
  wire [8:0] current_output = reg_[17:9]; // @[\\src\\main\\scala\\LFSR.scala 19:27]
  reg [9:0] history_0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_1; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_2; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_3; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_4; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_5; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_6; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_7; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_8; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_9; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_10; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_11; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_12; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_13; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_14; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_15; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_16; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_17; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_18; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_19; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_20; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_21; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_22; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_23; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_24; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_25; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_26; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_27; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_28; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_29; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  assign io_out_0 = history_0; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_1 = history_1; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_2 = history_2; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_3 = history_3; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_4 = history_4; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_5 = history_5; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_6 = history_6; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_7 = history_7; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_8 = history_8; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_9 = history_9; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_20 = history_20; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_21 = history_21; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_22 = history_22; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_23 = history_23; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_24 = history_24; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_25 = history_25; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_26 = history_26; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_27 = history_27; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_28 = history_28; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_29 = history_29; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 10:20]
      reg_ <= 64'h123456789abcdef; // @[\\src\\main\\scala\\LFSR.scala 10:20]
    end else begin
      reg_ <= _reg_T_1; // @[\\src\\main\\scala\\LFSR.scala 16:7]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_0 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_0 <= history_1; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_1 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_1 <= history_2; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_2 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_2 <= history_3; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_3 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_3 <= history_4; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_4 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_4 <= history_5; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_5 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_5 <= history_6; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_6 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_6 <= history_7; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_7 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_7 <= history_8; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_8 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_8 <= history_9; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_9 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_9 <= history_10; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_10 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_10 <= history_11; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_11 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_11 <= history_12; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_12 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_12 <= history_13; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_13 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_13 <= history_14; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_14 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_14 <= history_15; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_15 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_15 <= history_16; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_16 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_16 <= history_17; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_17 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_17 <= history_18; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_18 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_18 <= history_19; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_19 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_19 <= history_20; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_20 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_20 <= history_21; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_21 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_21 <= history_22; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_22 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_22 <= history_23; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_23 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_23 <= history_24; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_24 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_24 <= history_25; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_25 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_25 <= history_26; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_26 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_26 <= history_27; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_27 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_27 <= history_28; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_28 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_28 <= history_29; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_29 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_29 <= {{1'd0}, current_output}; // @[\\src\\main\\scala\\LFSR.scala 28:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_ = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  history_0 = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  history_1 = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  history_2 = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  history_3 = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  history_4 = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  history_5 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  history_6 = _RAND_7[9:0];
  _RAND_8 = {1{`RANDOM}};
  history_7 = _RAND_8[9:0];
  _RAND_9 = {1{`RANDOM}};
  history_8 = _RAND_9[9:0];
  _RAND_10 = {1{`RANDOM}};
  history_9 = _RAND_10[9:0];
  _RAND_11 = {1{`RANDOM}};
  history_10 = _RAND_11[9:0];
  _RAND_12 = {1{`RANDOM}};
  history_11 = _RAND_12[9:0];
  _RAND_13 = {1{`RANDOM}};
  history_12 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  history_13 = _RAND_14[9:0];
  _RAND_15 = {1{`RANDOM}};
  history_14 = _RAND_15[9:0];
  _RAND_16 = {1{`RANDOM}};
  history_15 = _RAND_16[9:0];
  _RAND_17 = {1{`RANDOM}};
  history_16 = _RAND_17[9:0];
  _RAND_18 = {1{`RANDOM}};
  history_17 = _RAND_18[9:0];
  _RAND_19 = {1{`RANDOM}};
  history_18 = _RAND_19[9:0];
  _RAND_20 = {1{`RANDOM}};
  history_19 = _RAND_20[9:0];
  _RAND_21 = {1{`RANDOM}};
  history_20 = _RAND_21[9:0];
  _RAND_22 = {1{`RANDOM}};
  history_21 = _RAND_22[9:0];
  _RAND_23 = {1{`RANDOM}};
  history_22 = _RAND_23[9:0];
  _RAND_24 = {1{`RANDOM}};
  history_23 = _RAND_24[9:0];
  _RAND_25 = {1{`RANDOM}};
  history_24 = _RAND_25[9:0];
  _RAND_26 = {1{`RANDOM}};
  history_25 = _RAND_26[9:0];
  _RAND_27 = {1{`RANDOM}};
  history_26 = _RAND_27[9:0];
  _RAND_28 = {1{`RANDOM}};
  history_27 = _RAND_28[9:0];
  _RAND_29 = {1{`RANDOM}};
  history_28 = _RAND_29[9:0];
  _RAND_30 = {1{`RANDOM}};
  history_29 = _RAND_30[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GameLogic(
  input         clock,
  input         reset,
  input         io_btnC, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnU, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnL, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnR, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnD, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_3, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_7, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_8, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_9, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_10, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_11, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_12, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_13, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_14, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_46, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_47, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_48, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_49, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_50, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_51, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_52, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_53, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_54, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_55, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_56, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_57, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_61, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_62, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_63, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_3, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_7, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_8, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_9, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_10, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_11, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_12, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_13, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_14, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_46, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_47, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_48, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_49, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_50, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_51, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_52, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_53, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_54, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_55, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_56, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_57, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_61, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_62, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_63, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_3, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_4, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_5, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_6, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_7, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_8, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_9, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_10, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_11, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_12, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_13, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_14, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_15, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_46, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_47, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_48, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_49, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_50, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_51, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_52, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_53, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_54, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_55, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_56, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_57, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_61, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_62, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_63, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_viewBoxX, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [8:0]  io_viewBoxY, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_newFrame, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_frameUpdateDone // @[\\src\\main\\scala\\GameLogic.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
`endif // RANDOMIZE_REG_INIT
  wire  difficulty_clock; // @[\\src\\main\\scala\\GameLogic.scala 210:26]
  wire  difficulty_reset; // @[\\src\\main\\scala\\GameLogic.scala 210:26]
  wire [1:0] difficulty_io_level; // @[\\src\\main\\scala\\GameLogic.scala 210:26]
  wire [26:0] difficulty_io_speed; // @[\\src\\main\\scala\\GameLogic.scala 210:26]
  wire  difficulty_io_resetSpeed; // @[\\src\\main\\scala\\GameLogic.scala 210:26]
  wire  lfsr_clock; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire  lfsr_reset; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_0; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_1; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_2; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_3; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_4; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_5; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_6; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_7; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_8; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_9; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_20; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_21; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_22; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_23; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_24; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_25; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_26; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_27; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_28; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  wire [9:0] lfsr_io_out_29; // @[\\src\\main\\scala\\GameLogic.scala 248:20]
  reg [2:0] stateReg; // @[\\src\\main\\scala\\GameLogic.scala 113:25]
  reg [10:0] spriteXRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [9:0] spriteYRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg  spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  initializePositions; // @[\\src\\main\\scala\\GameLogic.scala 131:36]
  wire [10:0] _GEN_0 = initializePositions ? $signed(11'sh140) : $signed(spriteXRegs_3); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_1 = initializePositions ? $signed(10'shf0) : $signed(spriteYRegs_3); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_14 = initializePositions ? $signed(11'sh140) : $signed(spriteXRegs_13); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_15 = initializePositions ? $signed(10'shf0) : $signed(spriteYRegs_13); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_16 = initializePositions ? $signed(11'sh260) : $signed(spriteXRegs_14); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_17 = initializePositions ? $signed(10'shf0) : $signed(spriteYRegs_14); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_18 = initializePositions ? $signed(11'sh168) : $signed(spriteXRegs_16); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_19 = initializePositions ? $signed(10'sh14) : $signed(spriteYRegs_16); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_20 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_17); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_21 = initializePositions ? $signed(10'sh32) : $signed(spriteYRegs_17); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_22 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_18); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_23 = initializePositions ? $signed(10'sh50) : $signed(spriteYRegs_18); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_24 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_19); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_25 = initializePositions ? $signed(10'sh6e) : $signed(spriteYRegs_19); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_26 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_20); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_27 = initializePositions ? $signed(10'sh8c) : $signed(spriteYRegs_20); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_28 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_21); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_29 = initializePositions ? $signed(10'shaa) : $signed(spriteYRegs_21); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_30 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_22); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_31 = initializePositions ? $signed(10'shc8) : $signed(spriteYRegs_22); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_32 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_23); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_33 = initializePositions ? $signed(10'she6) : $signed(spriteYRegs_23); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_34 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_24); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_35 = initializePositions ? $signed(10'sh104) : $signed(spriteYRegs_24); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_36 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_25); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_37 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_25); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_38 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_26); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_39 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_26); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_40 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_27); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_41 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_27); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_42 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_28); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_43 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_28); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_44 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_29); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_45 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_29); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_46 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_30); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_47 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_30); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_48 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_31); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_49 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_31); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_50 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_32); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_51 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_32); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_52 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_33); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_53 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_33); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_54 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_34); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_55 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_34); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_56 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_35); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_57 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_35); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_58 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_36); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_59 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_36); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_60 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_37); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_61 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_37); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_62 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_38); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_63 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_38); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_64 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_39); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_65 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_39); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_66 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_40); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_67 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_40); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_68 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_41); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_69 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_41); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_70 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_42); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_71 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_42); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_72 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_43); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_73 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_43); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_74 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_44); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_75 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_44); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_76 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_45); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_77 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_45); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_102 = initializePositions ? $signed(11'sh140) : $signed(spriteXRegs_58); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_103 = initializePositions ? $signed(10'sh14) : $signed(spriteYRegs_58); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_104 = initializePositions ? $signed(11'sh1f4) : $signed(spriteXRegs_59); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_105 = initializePositions ? $signed(10'sh46) : $signed(spriteYRegs_59); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire [10:0] _GEN_106 = initializePositions ? $signed(11'sh96) : $signed(spriteXRegs_60); // @[\\src\\main\\scala\\GameLogic.scala 132:29 162:23 121:28]
  wire [9:0] _GEN_107 = initializePositions ? $signed(10'sh64) : $signed(spriteYRegs_60); // @[\\src\\main\\scala\\GameLogic.scala 132:29 163:23 122:28]
  wire  _GEN_114 = initializePositions ? 1'h0 : initializePositions; // @[\\src\\main\\scala\\GameLogic.scala 132:29 165:25 131:36]
  reg  sprite58ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 169:42]
  reg  sprite58ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 170:40]
  reg  sprite59ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 171:42]
  reg  sprite59ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 172:40]
  reg  sprite60ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 173:42]
  reg  sprite60ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 174:40]
  reg [9:0] viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 202:28]
  reg [8:0] viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 203:28]
  reg [1:0] lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 212:23]
  reg [2:0] livesReg; // @[\\src\\main\\scala\\GameLogic.scala 223:25]
  reg [9:0] extraLifeCnt; // @[\\src\\main\\scala\\GameLogic.scala 226:29]
  wire  _difficulty_io_resetSpeed_T_1 = livesReg == 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 229:62]
  reg [7:0] spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 232:34]
  reg [5:0] nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 233:34]
  reg [9:0] starCnt; // @[\\src\\main\\scala\\GameLogic.scala 236:24]
  reg  collisionDetected; // @[\\src\\main\\scala\\GameLogic.scala 239:34]
  reg [7:0] blinkCounter; // @[\\src\\main\\scala\\GameLogic.scala 240:29]
  reg [1:0] blinkTimes; // @[\\src\\main\\scala\\GameLogic.scala 241:27]
  reg  isBlinking; // @[\\src\\main\\scala\\GameLogic.scala 242:27]
  wire  _T = lvlReg != 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 251:15]
  wire  _T_2 = livesReg == 3'h2; // @[\\src\\main\\scala\\GameLogic.scala 256:25]
  wire  _T_3 = livesReg == 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 260:25]
  wire  _GEN_117 = livesReg == 3'h2 | _T_3; // @[\\src\\main\\scala\\GameLogic.scala 256:34 257:29]
  wire  _GEN_120 = _difficulty_io_resetSpeed_T_1 | _GEN_117; // @[\\src\\main\\scala\\GameLogic.scala 252:28 253:29]
  wire  _GEN_121 = _difficulty_io_resetSpeed_T_1 | _T_2; // @[\\src\\main\\scala\\GameLogic.scala 252:28 254:29]
  wire  _GEN_123 = lvlReg != 2'h0 & _GEN_120; // @[\\src\\main\\scala\\GameLogic.scala 251:24 270:27]
  wire  _GEN_124 = lvlReg != 2'h0 & _GEN_121; // @[\\src\\main\\scala\\GameLogic.scala 251:24 271:27]
  wire  _GEN_125 = lvlReg != 2'h0 & _difficulty_io_resetSpeed_T_1; // @[\\src\\main\\scala\\GameLogic.scala 251:24 272:27]
  wire [9:0] _spriteYRegs_16_T_2 = 10'h64 + lfsr_io_out_0; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_417 = {{16{spriteXRegs_16[10]}},spriteXRegs_16}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_16_T_2 = $signed(_GEN_417) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_127 = spriteVisibleRegs_16 ? $signed(_spriteXRegs_16_T_2) : $signed({{16{_GEN_18[10]}},_GEN_18}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_128 = $signed(spriteXRegs_16) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_127); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_129 = $signed(spriteXRegs_16) >= 11'sh280 ? $signed(_spriteYRegs_16_T_2) : $signed(_GEN_19); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_130 = $signed(spriteXRegs_16) >= 11'sh280 ? lfsr_io_out_0[8] : spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_131 = ~spriteScaleTypeRegs_0 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [9:0] _spriteYRegs_17_T_2 = 10'h64 + lfsr_io_out_1; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_418 = {{16{spriteXRegs_17[10]}},spriteXRegs_17}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_17_T_2 = $signed(_GEN_418) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_132 = spriteVisibleRegs_17 ? $signed(_spriteXRegs_17_T_2) : $signed({{16{_GEN_20[10]}},_GEN_20}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_133 = $signed(spriteXRegs_17) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_132); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_134 = $signed(spriteXRegs_17) >= 11'sh280 ? $signed(_spriteYRegs_17_T_2) : $signed(_GEN_21); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_135 = $signed(spriteXRegs_17) >= 11'sh280 ? lfsr_io_out_1[8] : spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_136 = ~spriteScaleTypeRegs_1 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [9:0] _spriteYRegs_18_T_2 = 10'h64 + lfsr_io_out_2; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_419 = {{16{spriteXRegs_18[10]}},spriteXRegs_18}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_18_T_2 = $signed(_GEN_419) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_137 = spriteVisibleRegs_18 ? $signed(_spriteXRegs_18_T_2) : $signed({{16{_GEN_22[10]}},_GEN_22}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_138 = $signed(spriteXRegs_18) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_137); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_139 = $signed(spriteXRegs_18) >= 11'sh280 ? $signed(_spriteYRegs_18_T_2) : $signed(_GEN_23); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_140 = $signed(spriteXRegs_18) >= 11'sh280 ? lfsr_io_out_2[8] : spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_141 = ~spriteScaleTypeRegs_2 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [9:0] _spriteYRegs_19_T_2 = 10'h64 + lfsr_io_out_3; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_475 = {{16{spriteXRegs_19[10]}},spriteXRegs_19}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_19_T_2 = $signed(_GEN_475) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_142 = spriteVisibleRegs_19 ? $signed(_spriteXRegs_19_T_2) : $signed({{16{_GEN_24[10]}},_GEN_24}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_143 = $signed(spriteXRegs_19) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_142); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_144 = $signed(spriteXRegs_19) >= 11'sh280 ? $signed(_spriteYRegs_19_T_2) : $signed(_GEN_25); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_145 = $signed(spriteXRegs_19) >= 11'sh280 ? lfsr_io_out_3[8] : spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_146 = ~spriteScaleTypeRegs_3 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [9:0] _spriteYRegs_20_T_2 = 10'h64 + lfsr_io_out_4; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_476 = {{16{spriteXRegs_20[10]}},spriteXRegs_20}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_20_T_2 = $signed(_GEN_476) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_147 = spriteVisibleRegs_20 ? $signed(_spriteXRegs_20_T_2) : $signed({{16{_GEN_26[10]}},_GEN_26}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_148 = $signed(spriteXRegs_20) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_147); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_149 = $signed(spriteXRegs_20) >= 11'sh280 ? $signed(_spriteYRegs_20_T_2) : $signed(_GEN_27); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_150 = $signed(spriteXRegs_20) >= 11'sh280 ? lfsr_io_out_4[8] : spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_151 = ~spriteScaleTypeRegs_4 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [9:0] _spriteYRegs_21_T_2 = 10'h64 + lfsr_io_out_5; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_477 = {{16{spriteXRegs_21[10]}},spriteXRegs_21}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_21_T_2 = $signed(_GEN_477) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_152 = spriteVisibleRegs_21 ? $signed(_spriteXRegs_21_T_2) : $signed({{16{_GEN_28[10]}},_GEN_28}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_153 = $signed(spriteXRegs_21) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_152); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_154 = $signed(spriteXRegs_21) >= 11'sh280 ? $signed(_spriteYRegs_21_T_2) : $signed(_GEN_29); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_155 = $signed(spriteXRegs_21) >= 11'sh280 ? lfsr_io_out_5[8] : spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_156 = ~spriteScaleTypeRegs_5 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [9:0] _spriteYRegs_22_T_2 = 10'h64 + lfsr_io_out_6; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_482 = {{16{spriteXRegs_22[10]}},spriteXRegs_22}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_22_T_2 = $signed(_GEN_482) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_157 = spriteVisibleRegs_22 ? $signed(_spriteXRegs_22_T_2) : $signed({{16{_GEN_30[10]}},_GEN_30}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_158 = $signed(spriteXRegs_22) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_157); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_159 = $signed(spriteXRegs_22) >= 11'sh280 ? $signed(_spriteYRegs_22_T_2) : $signed(_GEN_31); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_160 = $signed(spriteXRegs_22) >= 11'sh280 ? lfsr_io_out_6[8] : spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_161 = ~spriteScaleTypeRegs_6 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [9:0] _spriteYRegs_23_T_2 = 10'h64 + lfsr_io_out_7; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_483 = {{16{spriteXRegs_23[10]}},spriteXRegs_23}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_23_T_2 = $signed(_GEN_483) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_162 = spriteVisibleRegs_23 ? $signed(_spriteXRegs_23_T_2) : $signed({{16{_GEN_32[10]}},_GEN_32}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_163 = $signed(spriteXRegs_23) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_162); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_164 = $signed(spriteXRegs_23) >= 11'sh280 ? $signed(_spriteYRegs_23_T_2) : $signed(_GEN_33); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_165 = $signed(spriteXRegs_23) >= 11'sh280 ? lfsr_io_out_7[8] : spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_166 = ~spriteScaleTypeRegs_7 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [9:0] _spriteYRegs_24_T_2 = 10'h64 + lfsr_io_out_8; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_484 = {{16{spriteXRegs_24[10]}},spriteXRegs_24}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_24_T_2 = $signed(_GEN_484) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_167 = spriteVisibleRegs_24 ? $signed(_spriteXRegs_24_T_2) : $signed({{16{_GEN_34[10]}},_GEN_34}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_168 = $signed(spriteXRegs_24) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_167); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_169 = $signed(spriteXRegs_24) >= 11'sh280 ? $signed(_spriteYRegs_24_T_2) : $signed(_GEN_35); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_170 = $signed(spriteXRegs_24) >= 11'sh280 ? lfsr_io_out_8[8] : spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_171 = ~spriteScaleTypeRegs_8 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [9:0] _spriteYRegs_25_T_2 = 10'h64 + lfsr_io_out_9; // @[\\src\\main\\scala\\GameLogic.scala 302:63]
  wire [26:0] _GEN_540 = {{16{spriteXRegs_25[10]}},spriteXRegs_25}; // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _spriteXRegs_25_T_2 = $signed(_GEN_540) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 307:46]
  wire [26:0] _GEN_172 = spriteVisibleRegs_25 ? $signed(_spriteXRegs_25_T_2) : $signed({{16{_GEN_36[10]}},_GEN_36}); // @[\\src\\main\\scala\\GameLogic.scala 306:44 307:28]
  wire [26:0] _GEN_173 = $signed(spriteXRegs_25) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_172); // @[\\src\\main\\scala\\GameLogic.scala 300:41 301:28]
  wire [9:0] _GEN_174 = $signed(spriteXRegs_25) >= 11'sh280 ? $signed(_spriteYRegs_25_T_2) : $signed(_GEN_37); // @[\\src\\main\\scala\\GameLogic.scala 300:41 302:28]
  wire  _GEN_175 = $signed(spriteXRegs_25) >= 11'sh280 ? lfsr_io_out_9[8] : spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 126:36 300:41 304:40]
  wire  _GEN_176 = ~spriteScaleTypeRegs_9 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 311:52 312:43 315:43]
  wire [26:0] _GEN_541 = {{16{spriteXRegs_26[10]}},spriteXRegs_26}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_26_T_2 = $signed(_GEN_541) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_177 = spriteVisibleRegs_26 ? $signed(_spriteXRegs_26_T_2) : $signed({{16{_GEN_38[10]}},_GEN_38}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_178 = $signed(spriteXRegs_26) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_177); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_179 = $signed(spriteXRegs_26) >= 11'sh280 ? $signed(_spriteYRegs_16_T_2) : $signed(_GEN_39); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_180 = $signed(spriteXRegs_26) >= 11'sh280 ? lfsr_io_out_0[8] : _GEN_130; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [26:0] _GEN_542 = {{16{spriteXRegs_27[10]}},spriteXRegs_27}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_27_T_2 = $signed(_GEN_542) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_182 = spriteVisibleRegs_27 ? $signed(_spriteXRegs_27_T_2) : $signed({{16{_GEN_40[10]}},_GEN_40}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_183 = $signed(spriteXRegs_27) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_182); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_184 = $signed(spriteXRegs_27) >= 11'sh280 ? $signed(_spriteYRegs_17_T_2) : $signed(_GEN_41); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_185 = $signed(spriteXRegs_27) >= 11'sh280 ? lfsr_io_out_1[8] : _GEN_135; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [26:0] _GEN_548 = {{16{spriteXRegs_28[10]}},spriteXRegs_28}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_28_T_2 = $signed(_GEN_548) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_187 = spriteVisibleRegs_28 ? $signed(_spriteXRegs_28_T_2) : $signed({{16{_GEN_42[10]}},_GEN_42}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_188 = $signed(spriteXRegs_28) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_187); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_189 = $signed(spriteXRegs_28) >= 11'sh280 ? $signed(_spriteYRegs_18_T_2) : $signed(_GEN_43); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_190 = $signed(spriteXRegs_28) >= 11'sh280 ? lfsr_io_out_2[8] : _GEN_140; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [26:0] _GEN_549 = {{16{spriteXRegs_29[10]}},spriteXRegs_29}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_29_T_2 = $signed(_GEN_549) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_192 = spriteVisibleRegs_29 ? $signed(_spriteXRegs_29_T_2) : $signed({{16{_GEN_44[10]}},_GEN_44}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_193 = $signed(spriteXRegs_29) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_192); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_194 = $signed(spriteXRegs_29) >= 11'sh280 ? $signed(_spriteYRegs_19_T_2) : $signed(_GEN_45); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_195 = $signed(spriteXRegs_29) >= 11'sh280 ? lfsr_io_out_3[8] : _GEN_145; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [26:0] _GEN_550 = {{16{spriteXRegs_30[10]}},spriteXRegs_30}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_30_T_2 = $signed(_GEN_550) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_197 = spriteVisibleRegs_30 ? $signed(_spriteXRegs_30_T_2) : $signed({{16{_GEN_46[10]}},_GEN_46}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_198 = $signed(spriteXRegs_30) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_197); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_199 = $signed(spriteXRegs_30) >= 11'sh280 ? $signed(_spriteYRegs_20_T_2) : $signed(_GEN_47); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_200 = $signed(spriteXRegs_30) >= 11'sh280 ? lfsr_io_out_4[8] : _GEN_150; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [26:0] _GEN_606 = {{16{spriteXRegs_31[10]}},spriteXRegs_31}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_31_T_2 = $signed(_GEN_606) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_202 = spriteVisibleRegs_31 ? $signed(_spriteXRegs_31_T_2) : $signed({{16{_GEN_48[10]}},_GEN_48}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_203 = $signed(spriteXRegs_31) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_202); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_204 = $signed(spriteXRegs_31) >= 11'sh280 ? $signed(_spriteYRegs_21_T_2) : $signed(_GEN_49); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_205 = $signed(spriteXRegs_31) >= 11'sh280 ? lfsr_io_out_5[8] : _GEN_155; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [26:0] _GEN_607 = {{16{spriteXRegs_32[10]}},spriteXRegs_32}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_32_T_2 = $signed(_GEN_607) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_207 = spriteVisibleRegs_32 ? $signed(_spriteXRegs_32_T_2) : $signed({{16{_GEN_50[10]}},_GEN_50}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_208 = $signed(spriteXRegs_32) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_207); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_209 = $signed(spriteXRegs_32) >= 11'sh280 ? $signed(_spriteYRegs_22_T_2) : $signed(_GEN_51); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_210 = $signed(spriteXRegs_32) >= 11'sh280 ? lfsr_io_out_6[8] : _GEN_160; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [26:0] _GEN_608 = {{16{spriteXRegs_33[10]}},spriteXRegs_33}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_33_T_2 = $signed(_GEN_608) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_212 = spriteVisibleRegs_33 ? $signed(_spriteXRegs_33_T_2) : $signed({{16{_GEN_52[10]}},_GEN_52}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_213 = $signed(spriteXRegs_33) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_212); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_214 = $signed(spriteXRegs_33) >= 11'sh280 ? $signed(_spriteYRegs_23_T_2) : $signed(_GEN_53); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_215 = $signed(spriteXRegs_33) >= 11'sh280 ? lfsr_io_out_7[8] : _GEN_165; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [26:0] _GEN_613 = {{16{spriteXRegs_34[10]}},spriteXRegs_34}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_34_T_2 = $signed(_GEN_613) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_217 = spriteVisibleRegs_34 ? $signed(_spriteXRegs_34_T_2) : $signed({{16{_GEN_54[10]}},_GEN_54}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_218 = $signed(spriteXRegs_34) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_217); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_219 = $signed(spriteXRegs_34) >= 11'sh280 ? $signed(_spriteYRegs_24_T_2) : $signed(_GEN_55); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_220 = $signed(spriteXRegs_34) >= 11'sh280 ? lfsr_io_out_8[8] : _GEN_170; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [26:0] _GEN_614 = {{16{spriteXRegs_35[10]}},spriteXRegs_35}; // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _spriteXRegs_35_T_2 = $signed(_GEN_614) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 330:46]
  wire [26:0] _GEN_222 = spriteVisibleRegs_35 ? $signed(_spriteXRegs_35_T_2) : $signed({{16{_GEN_56[10]}},_GEN_56}); // @[\\src\\main\\scala\\GameLogic.scala 329:44 330:28]
  wire [26:0] _GEN_223 = $signed(spriteXRegs_35) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_222); // @[\\src\\main\\scala\\GameLogic.scala 323:41 324:28]
  wire [9:0] _GEN_224 = $signed(spriteXRegs_35) >= 11'sh280 ? $signed(_spriteYRegs_25_T_2) : $signed(_GEN_57); // @[\\src\\main\\scala\\GameLogic.scala 323:41 325:28]
  wire  _GEN_225 = $signed(spriteXRegs_35) >= 11'sh280 ? lfsr_io_out_9[8] : _GEN_175; // @[\\src\\main\\scala\\GameLogic.scala 323:41 327:40]
  wire [9:0] _spriteYRegs_36_T_2 = 10'h64 + lfsr_io_out_20; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_615 = {{16{spriteXRegs_36[10]}},spriteXRegs_36}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_36_T_2 = $signed(_GEN_615) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_227 = spriteVisibleRegs_36 ? $signed(_spriteXRegs_36_T_2) : $signed({{16{_GEN_58[10]}},_GEN_58}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_228 = $signed(spriteXRegs_36) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_227); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_229 = $signed(spriteXRegs_36) >= 11'sh280 ? $signed(_spriteYRegs_36_T_2) : $signed(_GEN_59); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_230 = $signed(spriteXRegs_36) >= 11'sh280 ? lfsr_io_out_0[8] : _GEN_180; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _spriteYRegs_37_T_2 = 10'h64 + lfsr_io_out_21; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_671 = {{16{spriteXRegs_37[10]}},spriteXRegs_37}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_37_T_2 = $signed(_GEN_671) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_232 = spriteVisibleRegs_37 ? $signed(_spriteXRegs_37_T_2) : $signed({{16{_GEN_60[10]}},_GEN_60}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_233 = $signed(spriteXRegs_37) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_232); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_234 = $signed(spriteXRegs_37) >= 11'sh280 ? $signed(_spriteYRegs_37_T_2) : $signed(_GEN_61); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_235 = $signed(spriteXRegs_37) >= 11'sh280 ? lfsr_io_out_1[8] : _GEN_185; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _spriteYRegs_38_T_2 = 10'h64 + lfsr_io_out_22; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_672 = {{16{spriteXRegs_38[10]}},spriteXRegs_38}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_38_T_2 = $signed(_GEN_672) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_237 = spriteVisibleRegs_38 ? $signed(_spriteXRegs_38_T_2) : $signed({{16{_GEN_62[10]}},_GEN_62}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_238 = $signed(spriteXRegs_38) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_237); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_239 = $signed(spriteXRegs_38) >= 11'sh280 ? $signed(_spriteYRegs_38_T_2) : $signed(_GEN_63); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_240 = $signed(spriteXRegs_38) >= 11'sh280 ? lfsr_io_out_2[8] : _GEN_190; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _spriteYRegs_39_T_2 = 10'h64 + lfsr_io_out_23; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_673 = {{16{spriteXRegs_39[10]}},spriteXRegs_39}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_39_T_2 = $signed(_GEN_673) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_242 = spriteVisibleRegs_39 ? $signed(_spriteXRegs_39_T_2) : $signed({{16{_GEN_64[10]}},_GEN_64}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_243 = $signed(spriteXRegs_39) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_242); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_244 = $signed(spriteXRegs_39) >= 11'sh280 ? $signed(_spriteYRegs_39_T_2) : $signed(_GEN_65); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_245 = $signed(spriteXRegs_39) >= 11'sh280 ? lfsr_io_out_3[8] : _GEN_195; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _spriteYRegs_40_T_2 = 10'h64 + lfsr_io_out_24; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_679 = {{16{spriteXRegs_40[10]}},spriteXRegs_40}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_40_T_2 = $signed(_GEN_679) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_247 = spriteVisibleRegs_40 ? $signed(_spriteXRegs_40_T_2) : $signed({{16{_GEN_66[10]}},_GEN_66}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_248 = $signed(spriteXRegs_40) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_247); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_249 = $signed(spriteXRegs_40) >= 11'sh280 ? $signed(_spriteYRegs_40_T_2) : $signed(_GEN_67); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_250 = $signed(spriteXRegs_40) >= 11'sh280 ? lfsr_io_out_4[8] : _GEN_200; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _spriteYRegs_41_T_2 = 10'h64 + lfsr_io_out_25; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_680 = {{16{spriteXRegs_41[10]}},spriteXRegs_41}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_41_T_2 = $signed(_GEN_680) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_252 = spriteVisibleRegs_41 ? $signed(_spriteXRegs_41_T_2) : $signed({{16{_GEN_68[10]}},_GEN_68}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_253 = $signed(spriteXRegs_41) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_252); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_254 = $signed(spriteXRegs_41) >= 11'sh280 ? $signed(_spriteYRegs_41_T_2) : $signed(_GEN_69); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_255 = $signed(spriteXRegs_41) >= 11'sh280 ? lfsr_io_out_5[8] : _GEN_205; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _spriteYRegs_42_T_2 = 10'h64 + lfsr_io_out_26; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_681 = {{16{spriteXRegs_42[10]}},spriteXRegs_42}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_42_T_2 = $signed(_GEN_681) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_257 = spriteVisibleRegs_42 ? $signed(_spriteXRegs_42_T_2) : $signed({{16{_GEN_70[10]}},_GEN_70}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_258 = $signed(spriteXRegs_42) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_257); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_259 = $signed(spriteXRegs_42) >= 11'sh280 ? $signed(_spriteYRegs_42_T_2) : $signed(_GEN_71); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_260 = $signed(spriteXRegs_42) >= 11'sh280 ? lfsr_io_out_6[8] : _GEN_210; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _spriteYRegs_43_T_2 = 10'h64 + lfsr_io_out_27; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_737 = {{16{spriteXRegs_43[10]}},spriteXRegs_43}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_43_T_2 = $signed(_GEN_737) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_262 = spriteVisibleRegs_43 ? $signed(_spriteXRegs_43_T_2) : $signed({{16{_GEN_72[10]}},_GEN_72}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_263 = $signed(spriteXRegs_43) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_262); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_264 = $signed(spriteXRegs_43) >= 11'sh280 ? $signed(_spriteYRegs_43_T_2) : $signed(_GEN_73); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_265 = $signed(spriteXRegs_43) >= 11'sh280 ? lfsr_io_out_7[8] : _GEN_215; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _spriteYRegs_44_T_2 = 10'h64 + lfsr_io_out_28; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_738 = {{16{spriteXRegs_44[10]}},spriteXRegs_44}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_44_T_2 = $signed(_GEN_738) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_267 = spriteVisibleRegs_44 ? $signed(_spriteXRegs_44_T_2) : $signed({{16{_GEN_74[10]}},_GEN_74}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_268 = $signed(spriteXRegs_44) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_267); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_269 = $signed(spriteXRegs_44) >= 11'sh280 ? $signed(_spriteYRegs_44_T_2) : $signed(_GEN_75); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_270 = $signed(spriteXRegs_44) >= 11'sh280 ? lfsr_io_out_8[8] : _GEN_220; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _spriteYRegs_45_T_2 = 10'h64 + lfsr_io_out_29; // @[\\src\\main\\scala\\GameLogic.scala 348:63]
  wire [26:0] _GEN_739 = {{16{spriteXRegs_45[10]}},spriteXRegs_45}; // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _spriteXRegs_45_T_2 = $signed(_GEN_739) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 354:46]
  wire [26:0] _GEN_272 = spriteVisibleRegs_45 ? $signed(_spriteXRegs_45_T_2) : $signed({{16{_GEN_76[10]}},_GEN_76}); // @[\\src\\main\\scala\\GameLogic.scala 353:44 354:28]
  wire [26:0] _GEN_273 = $signed(spriteXRegs_45) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_272); // @[\\src\\main\\scala\\GameLogic.scala 346:41 347:28]
  wire [9:0] _GEN_274 = $signed(spriteXRegs_45) >= 11'sh280 ? $signed(_spriteYRegs_45_T_2) : $signed(_GEN_77); // @[\\src\\main\\scala\\GameLogic.scala 346:41 348:28]
  wire  _GEN_275 = $signed(spriteXRegs_45) >= 11'sh280 ? lfsr_io_out_9[8] : _GEN_225; // @[\\src\\main\\scala\\GameLogic.scala 346:41 351:40]
  wire [9:0] _extraLifeCnt_T_1 = extraLifeCnt + 10'h1; // @[\\src\\main\\scala\\GameLogic.scala 374:40]
  wire [10:0] _GEN_277 = extraLifeCnt == 10'h258 ? $signed(-11'sh20) : $signed(_GEN_14); // @[\\src\\main\\scala\\GameLogic.scala 368:38 369:27]
  wire  _GEN_278 = extraLifeCnt == 10'h258 | spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 368:38 370:33 125:34]
  wire [9:0] _GEN_279 = extraLifeCnt == 10'h258 ? $signed(lfsr_io_out_0) : $signed(_GEN_15); // @[\\src\\main\\scala\\GameLogic.scala 368:38 371:27]
  wire [9:0] _GEN_280 = extraLifeCnt == 10'h258 ? 10'h0 : _extraLifeCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 368:38 372:24 374:24]
  wire [10:0] _spriteXRegs_13_T_2 = $signed(spriteXRegs_13) + 11'sh2; // @[\\src\\main\\scala\\GameLogic.scala 377:46]
  wire [10:0] _GEN_281 = spriteVisibleRegs_13 ? $signed(_spriteXRegs_13_T_2) : $signed(_GEN_277); // @[\\src\\main\\scala\\GameLogic.scala 376:37 377:27]
  wire  _GEN_282 = $signed(spriteXRegs_13) >= 11'sh280 ? 1'h0 : _GEN_278; // @[\\src\\main\\scala\\GameLogic.scala 379:40 380:33]
  wire [26:0] _GEN_283 = _T ? $signed(_GEN_128) : $signed({{16{_GEN_18[10]}},_GEN_18}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_286 = _T ? _GEN_131 : spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_288 = _T ? $signed(_GEN_133) : $signed({{16{_GEN_20[10]}},_GEN_20}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_291 = _T ? _GEN_136 : spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_293 = _T ? $signed(_GEN_138) : $signed({{16{_GEN_22[10]}},_GEN_22}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_296 = _T ? _GEN_141 : spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_298 = _T ? $signed(_GEN_143) : $signed({{16{_GEN_24[10]}},_GEN_24}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_301 = _T ? _GEN_146 : spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_303 = _T ? $signed(_GEN_148) : $signed({{16{_GEN_26[10]}},_GEN_26}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_306 = _T ? _GEN_151 : spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_308 = _T ? $signed(_GEN_153) : $signed({{16{_GEN_28[10]}},_GEN_28}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_311 = _T ? _GEN_156 : spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_313 = _T ? $signed(_GEN_158) : $signed({{16{_GEN_30[10]}},_GEN_30}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_316 = _T ? _GEN_161 : spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_318 = _T ? $signed(_GEN_163) : $signed({{16{_GEN_32[10]}},_GEN_32}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_321 = _T ? _GEN_166 : spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_323 = _T ? $signed(_GEN_168) : $signed({{16{_GEN_34[10]}},_GEN_34}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_326 = _T ? _GEN_171 : spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_328 = _T ? $signed(_GEN_173) : $signed({{16{_GEN_36[10]}},_GEN_36}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_331 = _T ? _GEN_176 : spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 294:29 188:33]
  wire [26:0] _GEN_333 = _T ? $signed(_GEN_178) : $signed({{16{_GEN_38[10]}},_GEN_38}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_337 = _T ? $signed(_GEN_183) : $signed({{16{_GEN_40[10]}},_GEN_40}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_341 = _T ? $signed(_GEN_188) : $signed({{16{_GEN_42[10]}},_GEN_42}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_345 = _T ? $signed(_GEN_193) : $signed({{16{_GEN_44[10]}},_GEN_44}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_349 = _T ? $signed(_GEN_198) : $signed({{16{_GEN_46[10]}},_GEN_46}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_353 = _T ? $signed(_GEN_203) : $signed({{16{_GEN_48[10]}},_GEN_48}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_357 = _T ? $signed(_GEN_208) : $signed({{16{_GEN_50[10]}},_GEN_50}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_361 = _T ? $signed(_GEN_213) : $signed({{16{_GEN_52[10]}},_GEN_52}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_365 = _T ? $signed(_GEN_218) : $signed({{16{_GEN_54[10]}},_GEN_54}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_369 = _T ? $signed(_GEN_223) : $signed({{16{_GEN_56[10]}},_GEN_56}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_373 = _T ? $signed(_GEN_228) : $signed({{16{_GEN_58[10]}},_GEN_58}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_377 = _T ? $signed(_GEN_233) : $signed({{16{_GEN_60[10]}},_GEN_60}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_381 = _T ? $signed(_GEN_238) : $signed({{16{_GEN_62[10]}},_GEN_62}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_385 = _T ? $signed(_GEN_243) : $signed({{16{_GEN_64[10]}},_GEN_64}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_389 = _T ? $signed(_GEN_248) : $signed({{16{_GEN_66[10]}},_GEN_66}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_393 = _T ? $signed(_GEN_253) : $signed({{16{_GEN_68[10]}},_GEN_68}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_397 = _T ? $signed(_GEN_258) : $signed({{16{_GEN_70[10]}},_GEN_70}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_401 = _T ? $signed(_GEN_263) : $signed({{16{_GEN_72[10]}},_GEN_72}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_405 = _T ? $signed(_GEN_268) : $signed({{16{_GEN_74[10]}},_GEN_74}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire [26:0] _GEN_409 = _T ? $signed(_GEN_273) : $signed({{16{_GEN_76[10]}},_GEN_76}); // @[\\src\\main\\scala\\GameLogic.scala 294:29]
  wire  _GEN_414 = _T ? _GEN_282 : spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 294:29 125:34]
  wire  _T_68 = lvlReg == 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 385:19]
  wire  _T_71 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha; // @[\\src\\main\\scala\\GameLogic.scala 387:40]
  wire [5:0] _T_73 = 6'h10 + nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 388:34]
  wire  _GEN_420 = 6'h3 == _T_73 | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_421 = 6'h4 == _T_73 | spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_422 = 6'h5 == _T_73 | spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_423 = 6'h6 == _T_73 | spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_424 = 6'h7 == _T_73 | spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_425 = 6'h8 == _T_73 | spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_426 = 6'h9 == _T_73 | spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_427 = 6'ha == _T_73 | spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_428 = 6'hb == _T_73 | spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_429 = 6'hc == _T_73 | spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_430 = 6'hd == _T_73 | _GEN_414; // @[\\src\\main\\scala\\GameLogic.scala 388:{55,55}]
  wire  _GEN_431 = 6'he == _T_73 | spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_432 = 6'hf == _T_73 | spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_433 = 6'h10 == _T_73 | spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_434 = 6'h11 == _T_73 | spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_435 = 6'h12 == _T_73 | spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_436 = 6'h13 == _T_73 | spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_437 = 6'h14 == _T_73 | spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_438 = 6'h15 == _T_73 | spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_439 = 6'h16 == _T_73 | spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_440 = 6'h17 == _T_73 | spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_441 = 6'h18 == _T_73 | spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_442 = 6'h19 == _T_73 | spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_443 = 6'h1a == _T_73 | spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_444 = 6'h1b == _T_73 | spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_445 = 6'h1c == _T_73 | spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_446 = 6'h1d == _T_73 | spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_447 = 6'h1e == _T_73 | spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_448 = 6'h1f == _T_73 | spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_449 = 6'h20 == _T_73 | spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_450 = 6'h21 == _T_73 | spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_451 = 6'h22 == _T_73 | spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_452 = 6'h23 == _T_73 | spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_453 = 6'h24 == _T_73 | spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_454 = 6'h25 == _T_73 | spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_455 = 6'h26 == _T_73 | spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_456 = 6'h27 == _T_73 | spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_457 = 6'h28 == _T_73 | spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_458 = 6'h29 == _T_73 | spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_459 = 6'h2a == _T_73 | spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_460 = 6'h2b == _T_73 | spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_461 = 6'h2c == _T_73 | spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_462 = 6'h2d == _T_73 | spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_463 = 6'h2e == _T_73 | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_464 = 6'h2f == _T_73 | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_465 = 6'h30 == _T_73 | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_466 = 6'h31 == _T_73 | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_467 = 6'h32 == _T_73 | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_468 = 6'h33 == _T_73 | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_469 = 6'h34 == _T_73 | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_470 = 6'h35 == _T_73 | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_471 = 6'h36 == _T_73 | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_472 = 6'h37 == _T_73 | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_473 = 6'h38 == _T_73 | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_474 = 6'h39 == _T_73 | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 388:{55,55}]
  wire  _GEN_478 = 6'h3d == _T_73 | _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 388:{55,55}]
  wire  _GEN_479 = 6'h3e == _T_73 | _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 388:{55,55}]
  wire  _GEN_480 = 6'h3f == _T_73 | _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 388:{55,55}]
  wire [5:0] _nextSpriteToSpawn_T_1 = nextSpriteToSpawn + 6'h1; // @[\\src\\main\\scala\\GameLogic.scala 389:50]
  wire [7:0] _spawnDelayCounter_T_1 = spawnDelayCounter - 8'h1; // @[\\src\\main\\scala\\GameLogic.scala 392:50]
  wire [7:0] _GEN_481 = spawnDelayCounter > 8'h0 ? _spawnDelayCounter_T_1 : spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 391:45 392:29 232:34]
  wire  _GEN_485 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_420 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_486 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_421 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_487 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_422 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_488 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_423 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_489 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_424 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_490 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_425 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_491 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_426 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_492 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_427 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_493 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_428 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_494 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_429 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_495 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_430 : _GEN_414; // @[\\src\\main\\scala\\GameLogic.scala 387:69]
  wire  _GEN_496 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_431 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_497 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_432 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_498 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_433 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_499 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_434 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_500 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_435 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_501 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_436 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_502 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_437 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_503 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_438 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_504 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_439 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_505 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_440 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_506 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_441 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_507 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_442 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_508 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_443 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_509 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_444 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_510 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_445 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_511 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_446 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_512 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_447 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_513 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_448 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_514 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_449 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_515 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_450 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_516 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_451 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_517 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_452 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_518 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_453 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_519 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_454 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_520 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_455 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_521 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_456 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_522 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_457 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_523 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_458 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_524 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_459 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_525 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_460 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_526 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_461 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_527 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_462 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_528 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_463 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_529 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_464 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_530 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_465 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_531 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_466 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_532 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_467 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_533 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_468 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_534 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_469 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_535 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_470 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_536 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_471 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_537 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_472 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_538 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_473 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_539 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_474 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 387:69]
  wire  _GEN_543 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_478 : _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 387:69]
  wire  _GEN_544 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_479 : _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 387:69]
  wire  _GEN_545 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_480 : _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 387:69]
  wire [5:0] _GEN_546 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _nextSpriteToSpawn_T_1 :
    nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 387:69 389:29 233:34]
  wire [7:0] _GEN_547 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? 8'h1e : _GEN_481; // @[\\src\\main\\scala\\GameLogic.scala 387:69 390:29]
  wire  _T_75 = lvlReg == 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 394:25]
  wire [5:0] _T_80 = 6'h1a + nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 397:34]
  wire  _GEN_551 = 6'h3 == _T_80 | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_552 = 6'h4 == _T_80 | spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_553 = 6'h5 == _T_80 | spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_554 = 6'h6 == _T_80 | spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_555 = 6'h7 == _T_80 | spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_556 = 6'h8 == _T_80 | spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_557 = 6'h9 == _T_80 | spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_558 = 6'ha == _T_80 | spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_559 = 6'hb == _T_80 | spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_560 = 6'hc == _T_80 | spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_561 = 6'hd == _T_80 | _GEN_414; // @[\\src\\main\\scala\\GameLogic.scala 397:{55,55}]
  wire  _GEN_562 = 6'he == _T_80 | spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_563 = 6'hf == _T_80 | spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_564 = 6'h10 == _T_80 | spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_565 = 6'h11 == _T_80 | spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_566 = 6'h12 == _T_80 | spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_567 = 6'h13 == _T_80 | spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_568 = 6'h14 == _T_80 | spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_569 = 6'h15 == _T_80 | spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_570 = 6'h16 == _T_80 | spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_571 = 6'h17 == _T_80 | spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_572 = 6'h18 == _T_80 | spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_573 = 6'h19 == _T_80 | spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_574 = 6'h1a == _T_80 | spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_575 = 6'h1b == _T_80 | spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_576 = 6'h1c == _T_80 | spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_577 = 6'h1d == _T_80 | spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_578 = 6'h1e == _T_80 | spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_579 = 6'h1f == _T_80 | spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_580 = 6'h20 == _T_80 | spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_581 = 6'h21 == _T_80 | spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_582 = 6'h22 == _T_80 | spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_583 = 6'h23 == _T_80 | spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_584 = 6'h24 == _T_80 | spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_585 = 6'h25 == _T_80 | spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_586 = 6'h26 == _T_80 | spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_587 = 6'h27 == _T_80 | spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_588 = 6'h28 == _T_80 | spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_589 = 6'h29 == _T_80 | spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_590 = 6'h2a == _T_80 | spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_591 = 6'h2b == _T_80 | spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_592 = 6'h2c == _T_80 | spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_593 = 6'h2d == _T_80 | spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_594 = 6'h2e == _T_80 | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_595 = 6'h2f == _T_80 | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_596 = 6'h30 == _T_80 | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_597 = 6'h31 == _T_80 | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_598 = 6'h32 == _T_80 | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_599 = 6'h33 == _T_80 | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_600 = 6'h34 == _T_80 | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_601 = 6'h35 == _T_80 | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_602 = 6'h36 == _T_80 | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_603 = 6'h37 == _T_80 | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_604 = 6'h38 == _T_80 | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_605 = 6'h39 == _T_80 | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 397:{55,55}]
  wire  _GEN_609 = 6'h3d == _T_80 | _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 397:{55,55}]
  wire  _GEN_610 = 6'h3e == _T_80 | _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 397:{55,55}]
  wire  _GEN_611 = 6'h3f == _T_80 | _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 397:{55,55}]
  wire  _GEN_616 = _T_71 ? _GEN_551 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_617 = _T_71 ? _GEN_552 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_618 = _T_71 ? _GEN_553 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_619 = _T_71 ? _GEN_554 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_620 = _T_71 ? _GEN_555 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_621 = _T_71 ? _GEN_556 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_622 = _T_71 ? _GEN_557 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_623 = _T_71 ? _GEN_558 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_624 = _T_71 ? _GEN_559 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_625 = _T_71 ? _GEN_560 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_626 = _T_71 ? _GEN_561 : _GEN_414; // @[\\src\\main\\scala\\GameLogic.scala 396:69]
  wire  _GEN_627 = _T_71 ? _GEN_562 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_628 = _T_71 ? _GEN_563 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_629 = _T_71 ? _GEN_564 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_630 = _T_71 ? _GEN_565 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_631 = _T_71 ? _GEN_566 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_632 = _T_71 ? _GEN_567 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_633 = _T_71 ? _GEN_568 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_634 = _T_71 ? _GEN_569 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_635 = _T_71 ? _GEN_570 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_636 = _T_71 ? _GEN_571 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_637 = _T_71 ? _GEN_572 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_638 = _T_71 ? _GEN_573 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_639 = _T_71 ? _GEN_574 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_640 = _T_71 ? _GEN_575 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_641 = _T_71 ? _GEN_576 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_642 = _T_71 ? _GEN_577 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_643 = _T_71 ? _GEN_578 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_644 = _T_71 ? _GEN_579 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_645 = _T_71 ? _GEN_580 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_646 = _T_71 ? _GEN_581 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_647 = _T_71 ? _GEN_582 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_648 = _T_71 ? _GEN_583 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_649 = _T_71 ? _GEN_584 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_650 = _T_71 ? _GEN_585 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_651 = _T_71 ? _GEN_586 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_652 = _T_71 ? _GEN_587 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_653 = _T_71 ? _GEN_588 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_654 = _T_71 ? _GEN_589 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_655 = _T_71 ? _GEN_590 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_656 = _T_71 ? _GEN_591 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_657 = _T_71 ? _GEN_592 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_658 = _T_71 ? _GEN_593 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_659 = _T_71 ? _GEN_594 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_660 = _T_71 ? _GEN_595 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_661 = _T_71 ? _GEN_596 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_662 = _T_71 ? _GEN_597 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_663 = _T_71 ? _GEN_598 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_664 = _T_71 ? _GEN_599 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_665 = _T_71 ? _GEN_600 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_666 = _T_71 ? _GEN_601 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_667 = _T_71 ? _GEN_602 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_668 = _T_71 ? _GEN_603 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_669 = _T_71 ? _GEN_604 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_670 = _T_71 ? _GEN_605 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 396:69]
  wire  _GEN_674 = _T_71 ? _GEN_609 : _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 396:69]
  wire  _GEN_675 = _T_71 ? _GEN_610 : _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 396:69]
  wire  _GEN_676 = _T_71 ? _GEN_611 : _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 396:69]
  wire [7:0] _GEN_678 = _T_71 ? 8'h19 : _GEN_481; // @[\\src\\main\\scala\\GameLogic.scala 396:69 399:29]
  wire  _T_82 = lvlReg == 2'h3; // @[\\src\\main\\scala\\GameLogic.scala 403:25]
  wire [5:0] _T_87 = 6'h24 + nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 406:34]
  wire  _GEN_682 = 6'h3 == _T_87 | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_683 = 6'h4 == _T_87 | spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_684 = 6'h5 == _T_87 | spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_685 = 6'h6 == _T_87 | spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_686 = 6'h7 == _T_87 | spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_687 = 6'h8 == _T_87 | spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_688 = 6'h9 == _T_87 | spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_689 = 6'ha == _T_87 | spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_690 = 6'hb == _T_87 | spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_691 = 6'hc == _T_87 | spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_692 = 6'hd == _T_87 | _GEN_414; // @[\\src\\main\\scala\\GameLogic.scala 406:{55,55}]
  wire  _GEN_693 = 6'he == _T_87 | spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_694 = 6'hf == _T_87 | spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_695 = 6'h10 == _T_87 | spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_696 = 6'h11 == _T_87 | spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_697 = 6'h12 == _T_87 | spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_698 = 6'h13 == _T_87 | spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_699 = 6'h14 == _T_87 | spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_700 = 6'h15 == _T_87 | spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_701 = 6'h16 == _T_87 | spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_702 = 6'h17 == _T_87 | spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_703 = 6'h18 == _T_87 | spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_704 = 6'h19 == _T_87 | spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_705 = 6'h1a == _T_87 | spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_706 = 6'h1b == _T_87 | spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_707 = 6'h1c == _T_87 | spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_708 = 6'h1d == _T_87 | spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_709 = 6'h1e == _T_87 | spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_710 = 6'h1f == _T_87 | spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_711 = 6'h20 == _T_87 | spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_712 = 6'h21 == _T_87 | spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_713 = 6'h22 == _T_87 | spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_714 = 6'h23 == _T_87 | spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_715 = 6'h24 == _T_87 | spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_716 = 6'h25 == _T_87 | spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_717 = 6'h26 == _T_87 | spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_718 = 6'h27 == _T_87 | spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_719 = 6'h28 == _T_87 | spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_720 = 6'h29 == _T_87 | spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_721 = 6'h2a == _T_87 | spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_722 = 6'h2b == _T_87 | spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_723 = 6'h2c == _T_87 | spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_724 = 6'h2d == _T_87 | spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_725 = 6'h2e == _T_87 | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_726 = 6'h2f == _T_87 | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_727 = 6'h30 == _T_87 | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_728 = 6'h31 == _T_87 | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_729 = 6'h32 == _T_87 | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_730 = 6'h33 == _T_87 | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_731 = 6'h34 == _T_87 | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_732 = 6'h35 == _T_87 | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_733 = 6'h36 == _T_87 | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_734 = 6'h37 == _T_87 | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_735 = 6'h38 == _T_87 | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_736 = 6'h39 == _T_87 | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 406:{55,55}]
  wire  _GEN_740 = 6'h3d == _T_87 | _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 406:{55,55}]
  wire  _GEN_741 = 6'h3e == _T_87 | _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 406:{55,55}]
  wire  _GEN_742 = 6'h3f == _T_87 | _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 406:{55,55}]
  wire  _GEN_747 = _T_71 ? _GEN_682 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_748 = _T_71 ? _GEN_683 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_749 = _T_71 ? _GEN_684 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_750 = _T_71 ? _GEN_685 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_751 = _T_71 ? _GEN_686 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_752 = _T_71 ? _GEN_687 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_753 = _T_71 ? _GEN_688 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_754 = _T_71 ? _GEN_689 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_755 = _T_71 ? _GEN_690 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_756 = _T_71 ? _GEN_691 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_757 = _T_71 ? _GEN_692 : _GEN_414; // @[\\src\\main\\scala\\GameLogic.scala 405:69]
  wire  _GEN_758 = _T_71 ? _GEN_693 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_759 = _T_71 ? _GEN_694 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_760 = _T_71 ? _GEN_695 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_761 = _T_71 ? _GEN_696 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_762 = _T_71 ? _GEN_697 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_763 = _T_71 ? _GEN_698 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_764 = _T_71 ? _GEN_699 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_765 = _T_71 ? _GEN_700 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_766 = _T_71 ? _GEN_701 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_767 = _T_71 ? _GEN_702 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_768 = _T_71 ? _GEN_703 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_769 = _T_71 ? _GEN_704 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_770 = _T_71 ? _GEN_705 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_771 = _T_71 ? _GEN_706 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_772 = _T_71 ? _GEN_707 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_773 = _T_71 ? _GEN_708 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_774 = _T_71 ? _GEN_709 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_775 = _T_71 ? _GEN_710 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_776 = _T_71 ? _GEN_711 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_777 = _T_71 ? _GEN_712 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_778 = _T_71 ? _GEN_713 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_779 = _T_71 ? _GEN_714 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_780 = _T_71 ? _GEN_715 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_781 = _T_71 ? _GEN_716 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_782 = _T_71 ? _GEN_717 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_783 = _T_71 ? _GEN_718 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_784 = _T_71 ? _GEN_719 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_785 = _T_71 ? _GEN_720 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_786 = _T_71 ? _GEN_721 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_787 = _T_71 ? _GEN_722 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_788 = _T_71 ? _GEN_723 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_789 = _T_71 ? _GEN_724 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_790 = _T_71 ? _GEN_725 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_791 = _T_71 ? _GEN_726 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_792 = _T_71 ? _GEN_727 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_793 = _T_71 ? _GEN_728 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_794 = _T_71 ? _GEN_729 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_795 = _T_71 ? _GEN_730 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_796 = _T_71 ? _GEN_731 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_797 = _T_71 ? _GEN_732 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_798 = _T_71 ? _GEN_733 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_799 = _T_71 ? _GEN_734 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_800 = _T_71 ? _GEN_735 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_801 = _T_71 ? _GEN_736 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 405:69]
  wire  _GEN_805 = _T_71 ? _GEN_740 : _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 405:69]
  wire  _GEN_806 = _T_71 ? _GEN_741 : _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 405:69]
  wire  _GEN_807 = _T_71 ? _GEN_742 : _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 405:69]
  wire [7:0] _GEN_809 = _T_71 ? 8'h14 : _GEN_481; // @[\\src\\main\\scala\\GameLogic.scala 405:69 408:29]
  wire  _GEN_813 = lvlReg == 2'h3 ? _GEN_747 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_814 = lvlReg == 2'h3 ? _GEN_748 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_815 = lvlReg == 2'h3 ? _GEN_749 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_816 = lvlReg == 2'h3 ? _GEN_750 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_817 = lvlReg == 2'h3 ? _GEN_751 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_818 = lvlReg == 2'h3 ? _GEN_752 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_819 = lvlReg == 2'h3 ? _GEN_753 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_820 = lvlReg == 2'h3 ? _GEN_754 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_821 = lvlReg == 2'h3 ? _GEN_755 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_822 = lvlReg == 2'h3 ? _GEN_756 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_823 = lvlReg == 2'h3 ? _GEN_757 : _GEN_414; // @[\\src\\main\\scala\\GameLogic.scala 403:34]
  wire  _GEN_824 = lvlReg == 2'h3 ? _GEN_758 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_825 = lvlReg == 2'h3 ? _GEN_759 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_826 = lvlReg == 2'h3 ? _GEN_760 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_827 = lvlReg == 2'h3 ? _GEN_761 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_828 = lvlReg == 2'h3 ? _GEN_762 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_829 = lvlReg == 2'h3 ? _GEN_763 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_830 = lvlReg == 2'h3 ? _GEN_764 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_831 = lvlReg == 2'h3 ? _GEN_765 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_832 = lvlReg == 2'h3 ? _GEN_766 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_833 = lvlReg == 2'h3 ? _GEN_767 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_834 = lvlReg == 2'h3 ? _GEN_768 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_835 = lvlReg == 2'h3 ? _GEN_769 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_836 = lvlReg == 2'h3 ? _GEN_770 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_837 = lvlReg == 2'h3 ? _GEN_771 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_838 = lvlReg == 2'h3 ? _GEN_772 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_839 = lvlReg == 2'h3 ? _GEN_773 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_840 = lvlReg == 2'h3 ? _GEN_774 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_841 = lvlReg == 2'h3 ? _GEN_775 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_842 = lvlReg == 2'h3 ? _GEN_776 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_843 = lvlReg == 2'h3 ? _GEN_777 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_844 = lvlReg == 2'h3 ? _GEN_778 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_845 = lvlReg == 2'h3 ? _GEN_779 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_846 = lvlReg == 2'h3 ? _GEN_780 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_847 = lvlReg == 2'h3 ? _GEN_781 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_848 = lvlReg == 2'h3 ? _GEN_782 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_849 = lvlReg == 2'h3 ? _GEN_783 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_850 = lvlReg == 2'h3 ? _GEN_784 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_851 = lvlReg == 2'h3 ? _GEN_785 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_852 = lvlReg == 2'h3 ? _GEN_786 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_853 = lvlReg == 2'h3 ? _GEN_787 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_854 = lvlReg == 2'h3 ? _GEN_788 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_855 = lvlReg == 2'h3 ? _GEN_789 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_856 = lvlReg == 2'h3 ? _GEN_790 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_857 = lvlReg == 2'h3 ? _GEN_791 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_858 = lvlReg == 2'h3 ? _GEN_792 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_859 = lvlReg == 2'h3 ? _GEN_793 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_860 = lvlReg == 2'h3 ? _GEN_794 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_861 = lvlReg == 2'h3 ? _GEN_795 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_862 = lvlReg == 2'h3 ? _GEN_796 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_863 = lvlReg == 2'h3 ? _GEN_797 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_864 = lvlReg == 2'h3 ? _GEN_798 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_865 = lvlReg == 2'h3 ? _GEN_799 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_866 = lvlReg == 2'h3 ? _GEN_800 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_867 = lvlReg == 2'h3 ? _GEN_801 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 403:34]
  wire  _GEN_871 = lvlReg == 2'h3 ? _GEN_805 : _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 403:34]
  wire  _GEN_872 = lvlReg == 2'h3 ? _GEN_806 : _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 403:34]
  wire  _GEN_873 = lvlReg == 2'h3 ? _GEN_807 : _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 403:34]
  wire [5:0] _GEN_874 = lvlReg == 2'h3 ? _GEN_546 : nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 233:34 403:34]
  wire [7:0] _GEN_875 = lvlReg == 2'h3 ? _GEN_809 : spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 232:34 403:34]
  wire  _GEN_879 = lvlReg == 2'h2 ? _GEN_616 : _GEN_813; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_880 = lvlReg == 2'h2 ? _GEN_617 : _GEN_814; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_881 = lvlReg == 2'h2 ? _GEN_618 : _GEN_815; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_882 = lvlReg == 2'h2 ? _GEN_619 : _GEN_816; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_883 = lvlReg == 2'h2 ? _GEN_620 : _GEN_817; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_884 = lvlReg == 2'h2 ? _GEN_621 : _GEN_818; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_885 = lvlReg == 2'h2 ? _GEN_622 : _GEN_819; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_886 = lvlReg == 2'h2 ? _GEN_623 : _GEN_820; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_887 = lvlReg == 2'h2 ? _GEN_624 : _GEN_821; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_888 = lvlReg == 2'h2 ? _GEN_625 : _GEN_822; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_889 = lvlReg == 2'h2 ? _GEN_626 : _GEN_823; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_890 = lvlReg == 2'h2 ? _GEN_627 : _GEN_824; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_891 = lvlReg == 2'h2 ? _GEN_628 : _GEN_825; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_892 = lvlReg == 2'h2 ? _GEN_629 : _GEN_826; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_893 = lvlReg == 2'h2 ? _GEN_630 : _GEN_827; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_894 = lvlReg == 2'h2 ? _GEN_631 : _GEN_828; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_895 = lvlReg == 2'h2 ? _GEN_632 : _GEN_829; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_896 = lvlReg == 2'h2 ? _GEN_633 : _GEN_830; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_897 = lvlReg == 2'h2 ? _GEN_634 : _GEN_831; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_898 = lvlReg == 2'h2 ? _GEN_635 : _GEN_832; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_899 = lvlReg == 2'h2 ? _GEN_636 : _GEN_833; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_900 = lvlReg == 2'h2 ? _GEN_637 : _GEN_834; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_901 = lvlReg == 2'h2 ? _GEN_638 : _GEN_835; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_902 = lvlReg == 2'h2 ? _GEN_639 : _GEN_836; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_903 = lvlReg == 2'h2 ? _GEN_640 : _GEN_837; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_904 = lvlReg == 2'h2 ? _GEN_641 : _GEN_838; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_905 = lvlReg == 2'h2 ? _GEN_642 : _GEN_839; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_906 = lvlReg == 2'h2 ? _GEN_643 : _GEN_840; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_907 = lvlReg == 2'h2 ? _GEN_644 : _GEN_841; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_908 = lvlReg == 2'h2 ? _GEN_645 : _GEN_842; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_909 = lvlReg == 2'h2 ? _GEN_646 : _GEN_843; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_910 = lvlReg == 2'h2 ? _GEN_647 : _GEN_844; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_911 = lvlReg == 2'h2 ? _GEN_648 : _GEN_845; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_912 = lvlReg == 2'h2 ? _GEN_649 : _GEN_846; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_913 = lvlReg == 2'h2 ? _GEN_650 : _GEN_847; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_914 = lvlReg == 2'h2 ? _GEN_651 : _GEN_848; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_915 = lvlReg == 2'h2 ? _GEN_652 : _GEN_849; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_916 = lvlReg == 2'h2 ? _GEN_653 : _GEN_850; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_917 = lvlReg == 2'h2 ? _GEN_654 : _GEN_851; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_918 = lvlReg == 2'h2 ? _GEN_655 : _GEN_852; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_919 = lvlReg == 2'h2 ? _GEN_656 : _GEN_853; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_920 = lvlReg == 2'h2 ? _GEN_657 : _GEN_854; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_921 = lvlReg == 2'h2 ? _GEN_658 : _GEN_855; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_922 = lvlReg == 2'h2 ? _GEN_659 : _GEN_856; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_923 = lvlReg == 2'h2 ? _GEN_660 : _GEN_857; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_924 = lvlReg == 2'h2 ? _GEN_661 : _GEN_858; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_925 = lvlReg == 2'h2 ? _GEN_662 : _GEN_859; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_926 = lvlReg == 2'h2 ? _GEN_663 : _GEN_860; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_927 = lvlReg == 2'h2 ? _GEN_664 : _GEN_861; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_928 = lvlReg == 2'h2 ? _GEN_665 : _GEN_862; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_929 = lvlReg == 2'h2 ? _GEN_666 : _GEN_863; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_930 = lvlReg == 2'h2 ? _GEN_667 : _GEN_864; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_931 = lvlReg == 2'h2 ? _GEN_668 : _GEN_865; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_932 = lvlReg == 2'h2 ? _GEN_669 : _GEN_866; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_933 = lvlReg == 2'h2 ? _GEN_670 : _GEN_867; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_937 = lvlReg == 2'h2 ? _GEN_674 : _GEN_871; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_938 = lvlReg == 2'h2 ? _GEN_675 : _GEN_872; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_939 = lvlReg == 2'h2 ? _GEN_676 : _GEN_873; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire [5:0] _GEN_940 = lvlReg == 2'h2 ? _GEN_546 : _GEN_874; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire [7:0] _GEN_941 = lvlReg == 2'h2 ? _GEN_678 : _GEN_875; // @[\\src\\main\\scala\\GameLogic.scala 394:34]
  wire  _GEN_955 = lvlReg == 2'h1 ? _GEN_495 : _GEN_889; // @[\\src\\main\\scala\\GameLogic.scala 385:28]
  wire  _GEN_956 = lvlReg == 2'h1 ? _GEN_496 : _GEN_890; // @[\\src\\main\\scala\\GameLogic.scala 385:28]
  wire  _T_89 = ~isBlinking; // @[\\src\\main\\scala\\GameLogic.scala 417:12]
  wire [10:0] _T_94 = $signed(spriteXRegs_16) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_95 = $signed(spriteXRegs_14) < $signed(_T_94); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_96 = spriteVisibleRegs_16 & $signed(spriteXRegs_16) <= 11'sh280 & _T_95; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [10:0] _T_99 = $signed(spriteXRegs_14) + 11'sh8; // @[\\src\\main\\scala\\GameLogic.scala 421:94]
  wire [9:0] _T_104 = $signed(spriteYRegs_16) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_105 = $signed(spriteYRegs_14) < $signed(_T_104); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_106 = _T_96 & $signed(spriteXRegs_16) < $signed(_T_99) & _T_105; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire [9:0] _T_109 = $signed(spriteYRegs_14) + 10'shb; // @[\\src\\main\\scala\\GameLogic.scala 422:94]
  wire  _T_111 = _T_106 & $signed(spriteYRegs_16) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire  _GEN_1008 = _T_111 | collisionDetected; // @[\\src\\main\\scala\\GameLogic.scala 423:13 424:31 239:34]
  wire [10:0] _T_116 = $signed(spriteXRegs_17) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_117 = $signed(spriteXRegs_14) < $signed(_T_116); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_118 = spriteVisibleRegs_17 & $signed(spriteXRegs_17) <= 11'sh280 & _T_117; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [9:0] _T_126 = $signed(spriteYRegs_17) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_127 = $signed(spriteYRegs_14) < $signed(_T_126); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_128 = _T_118 & $signed(spriteXRegs_17) < $signed(_T_99) & _T_127; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire  _T_133 = _T_128 & $signed(spriteYRegs_17) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire [10:0] _T_138 = $signed(spriteXRegs_18) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_139 = $signed(spriteXRegs_14) < $signed(_T_138); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_140 = spriteVisibleRegs_18 & $signed(spriteXRegs_18) <= 11'sh280 & _T_139; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [9:0] _T_148 = $signed(spriteYRegs_18) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_149 = $signed(spriteYRegs_14) < $signed(_T_148); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_150 = _T_140 & $signed(spriteXRegs_18) < $signed(_T_99) & _T_149; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire  _T_155 = _T_150 & $signed(spriteYRegs_18) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire [10:0] _T_160 = $signed(spriteXRegs_19) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_161 = $signed(spriteXRegs_14) < $signed(_T_160); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_162 = spriteVisibleRegs_19 & $signed(spriteXRegs_19) <= 11'sh280 & _T_161; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [9:0] _T_170 = $signed(spriteYRegs_19) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_171 = $signed(spriteYRegs_14) < $signed(_T_170); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_172 = _T_162 & $signed(spriteXRegs_19) < $signed(_T_99) & _T_171; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire  _T_177 = _T_172 & $signed(spriteYRegs_19) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire [10:0] _T_182 = $signed(spriteXRegs_20) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_183 = $signed(spriteXRegs_14) < $signed(_T_182); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_184 = spriteVisibleRegs_20 & $signed(spriteXRegs_20) <= 11'sh280 & _T_183; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [9:0] _T_192 = $signed(spriteYRegs_20) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_193 = $signed(spriteYRegs_14) < $signed(_T_192); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_194 = _T_184 & $signed(spriteXRegs_20) < $signed(_T_99) & _T_193; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire  _T_199 = _T_194 & $signed(spriteYRegs_20) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire [10:0] _T_204 = $signed(spriteXRegs_21) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_205 = $signed(spriteXRegs_14) < $signed(_T_204); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_206 = spriteVisibleRegs_21 & $signed(spriteXRegs_21) <= 11'sh280 & _T_205; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [9:0] _T_214 = $signed(spriteYRegs_21) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_215 = $signed(spriteYRegs_14) < $signed(_T_214); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_216 = _T_206 & $signed(spriteXRegs_21) < $signed(_T_99) & _T_215; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire  _T_221 = _T_216 & $signed(spriteYRegs_21) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire [10:0] _T_226 = $signed(spriteXRegs_22) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_227 = $signed(spriteXRegs_14) < $signed(_T_226); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_228 = spriteVisibleRegs_22 & $signed(spriteXRegs_22) <= 11'sh280 & _T_227; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [9:0] _T_236 = $signed(spriteYRegs_22) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_237 = $signed(spriteYRegs_14) < $signed(_T_236); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_238 = _T_228 & $signed(spriteXRegs_22) < $signed(_T_99) & _T_237; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire  _T_243 = _T_238 & $signed(spriteYRegs_22) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire [10:0] _T_248 = $signed(spriteXRegs_23) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_249 = $signed(spriteXRegs_14) < $signed(_T_248); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_250 = spriteVisibleRegs_23 & $signed(spriteXRegs_23) <= 11'sh280 & _T_249; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [9:0] _T_258 = $signed(spriteYRegs_23) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_259 = $signed(spriteYRegs_14) < $signed(_T_258); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_260 = _T_250 & $signed(spriteXRegs_23) < $signed(_T_99) & _T_259; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire  _T_265 = _T_260 & $signed(spriteYRegs_23) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire [10:0] _T_270 = $signed(spriteXRegs_24) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_271 = $signed(spriteXRegs_14) < $signed(_T_270); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_272 = spriteVisibleRegs_24 & $signed(spriteXRegs_24) <= 11'sh280 & _T_271; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [9:0] _T_280 = $signed(spriteYRegs_24) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_281 = $signed(spriteYRegs_14) < $signed(_T_280); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_282 = _T_272 & $signed(spriteXRegs_24) < $signed(_T_99) & _T_281; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire  _T_287 = _T_282 & $signed(spriteYRegs_24) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire [10:0] _T_292 = $signed(spriteXRegs_25) + 11'sh1a; // @[\\src\\main\\scala\\GameLogic.scala 421:49]
  wire  _T_293 = $signed(spriteXRegs_14) < $signed(_T_292); // @[\\src\\main\\scala\\GameLogic.scala 421:32]
  wire  _T_294 = spriteVisibleRegs_25 & $signed(spriteXRegs_25) <= 11'sh280 & _T_293; // @[\\src\\main\\scala\\GameLogic.scala 420:63]
  wire [9:0] _T_302 = $signed(spriteYRegs_25) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 422:49]
  wire  _T_303 = $signed(spriteYRegs_14) < $signed(_T_302); // @[\\src\\main\\scala\\GameLogic.scala 422:32]
  wire  _T_304 = _T_294 & $signed(spriteXRegs_25) < $signed(_T_99) & _T_303; // @[\\src\\main\\scala\\GameLogic.scala 421:101]
  wire  _T_309 = _T_304 & $signed(spriteYRegs_25) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 422:57]
  wire  _GEN_1017 = _T_309 | (_T_287 | (_T_265 | (_T_243 | (_T_221 | (_T_199 | (_T_177 | (_T_155 | (_T_133 | _GEN_1008))
    )))))); // @[\\src\\main\\scala\\GameLogic.scala 423:13 424:31]
  wire  _GEN_1018 = ~isBlinking ? _GEN_1017 : collisionDetected; // @[\\src\\main\\scala\\GameLogic.scala 417:25 239:34]
  wire [10:0] _T_313 = $signed(spriteXRegs_26) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_314 = $signed(spriteXRegs_14) < $signed(_T_313); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_315 = spriteVisibleRegs_26 & _T_314; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_323 = $signed(spriteYRegs_26) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_324 = $signed(spriteYRegs_14) < $signed(_T_323); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_325 = _T_315 & $signed(spriteXRegs_26) < $signed(_T_99) & _T_324; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_330 = _T_325 & $signed(spriteYRegs_26) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire [10:0] _T_333 = $signed(spriteXRegs_27) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_334 = $signed(spriteXRegs_14) < $signed(_T_333); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_335 = spriteVisibleRegs_27 & _T_334; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_343 = $signed(spriteYRegs_27) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_344 = $signed(spriteYRegs_14) < $signed(_T_343); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_345 = _T_335 & $signed(spriteXRegs_27) < $signed(_T_99) & _T_344; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_350 = _T_345 & $signed(spriteYRegs_27) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire [10:0] _T_353 = $signed(spriteXRegs_28) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_354 = $signed(spriteXRegs_14) < $signed(_T_353); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_355 = spriteVisibleRegs_28 & _T_354; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_363 = $signed(spriteYRegs_28) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_364 = $signed(spriteYRegs_14) < $signed(_T_363); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_365 = _T_355 & $signed(spriteXRegs_28) < $signed(_T_99) & _T_364; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_370 = _T_365 & $signed(spriteYRegs_28) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire [10:0] _T_373 = $signed(spriteXRegs_29) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_374 = $signed(spriteXRegs_14) < $signed(_T_373); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_375 = spriteVisibleRegs_29 & _T_374; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_383 = $signed(spriteYRegs_29) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_384 = $signed(spriteYRegs_14) < $signed(_T_383); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_385 = _T_375 & $signed(spriteXRegs_29) < $signed(_T_99) & _T_384; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_390 = _T_385 & $signed(spriteYRegs_29) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire [10:0] _T_393 = $signed(spriteXRegs_30) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_394 = $signed(spriteXRegs_14) < $signed(_T_393); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_395 = spriteVisibleRegs_30 & _T_394; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_403 = $signed(spriteYRegs_30) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_404 = $signed(spriteYRegs_14) < $signed(_T_403); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_405 = _T_395 & $signed(spriteXRegs_30) < $signed(_T_99) & _T_404; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_410 = _T_405 & $signed(spriteYRegs_30) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire [10:0] _T_413 = $signed(spriteXRegs_31) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_414 = $signed(spriteXRegs_14) < $signed(_T_413); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_415 = spriteVisibleRegs_31 & _T_414; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_423 = $signed(spriteYRegs_31) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_424 = $signed(spriteYRegs_14) < $signed(_T_423); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_425 = _T_415 & $signed(spriteXRegs_31) < $signed(_T_99) & _T_424; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_430 = _T_425 & $signed(spriteYRegs_31) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire [10:0] _T_433 = $signed(spriteXRegs_32) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_434 = $signed(spriteXRegs_14) < $signed(_T_433); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_435 = spriteVisibleRegs_32 & _T_434; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_443 = $signed(spriteYRegs_32) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_444 = $signed(spriteYRegs_14) < $signed(_T_443); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_445 = _T_435 & $signed(spriteXRegs_32) < $signed(_T_99) & _T_444; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_450 = _T_445 & $signed(spriteYRegs_32) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire [10:0] _T_453 = $signed(spriteXRegs_33) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_454 = $signed(spriteXRegs_14) < $signed(_T_453); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_455 = spriteVisibleRegs_33 & _T_454; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_463 = $signed(spriteYRegs_33) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_464 = $signed(spriteYRegs_14) < $signed(_T_463); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_465 = _T_455 & $signed(spriteXRegs_33) < $signed(_T_99) & _T_464; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_470 = _T_465 & $signed(spriteYRegs_33) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire [10:0] _T_473 = $signed(spriteXRegs_34) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_474 = $signed(spriteXRegs_14) < $signed(_T_473); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_475 = spriteVisibleRegs_34 & _T_474; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_483 = $signed(spriteYRegs_34) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_484 = $signed(spriteYRegs_14) < $signed(_T_483); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_485 = _T_475 & $signed(spriteXRegs_34) < $signed(_T_99) & _T_484; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_490 = _T_485 & $signed(spriteYRegs_34) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire [10:0] _T_493 = $signed(spriteXRegs_35) + 11'sh1d; // @[\\src\\main\\scala\\GameLogic.scala 433:49]
  wire  _T_494 = $signed(spriteXRegs_14) < $signed(_T_493); // @[\\src\\main\\scala\\GameLogic.scala 433:32]
  wire  _T_495 = spriteVisibleRegs_35 & _T_494; // @[\\src\\main\\scala\\GameLogic.scala 432:34]
  wire [9:0] _T_503 = $signed(spriteYRegs_35) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 434:49]
  wire  _T_504 = $signed(spriteYRegs_14) < $signed(_T_503); // @[\\src\\main\\scala\\GameLogic.scala 434:32]
  wire  _T_505 = _T_495 & $signed(spriteXRegs_35) < $signed(_T_99) & _T_504; // @[\\src\\main\\scala\\GameLogic.scala 433:101]
  wire  _T_510 = _T_505 & $signed(spriteYRegs_35) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 434:57]
  wire  _GEN_1028 = _T_510 | (_T_490 | (_T_470 | (_T_450 | (_T_430 | (_T_410 | (_T_390 | (_T_370 | (_T_350 | (_T_330 |
    _GEN_1018))))))))); // @[\\src\\main\\scala\\GameLogic.scala 435:13 436:31]
  wire  _GEN_1029 = _T_89 ? _GEN_1028 : _GEN_1018; // @[\\src\\main\\scala\\GameLogic.scala 429:25]
  wire [10:0] _T_514 = $signed(spriteXRegs_36) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_515 = $signed(spriteXRegs_14) < $signed(_T_514); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_516 = spriteVisibleRegs_36 & _T_515; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_524 = $signed(spriteYRegs_36) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_525 = $signed(spriteYRegs_14) < $signed(_T_524); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_526 = _T_516 & $signed(spriteXRegs_36) < $signed(_T_99) & _T_525; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_531 = _T_526 & $signed(spriteYRegs_36) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire [10:0] _T_534 = $signed(spriteXRegs_37) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_535 = $signed(spriteXRegs_14) < $signed(_T_534); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_536 = spriteVisibleRegs_37 & _T_535; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_544 = $signed(spriteYRegs_37) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_545 = $signed(spriteYRegs_14) < $signed(_T_544); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_546 = _T_536 & $signed(spriteXRegs_37) < $signed(_T_99) & _T_545; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_551 = _T_546 & $signed(spriteYRegs_37) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire [10:0] _T_554 = $signed(spriteXRegs_38) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_555 = $signed(spriteXRegs_14) < $signed(_T_554); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_556 = spriteVisibleRegs_38 & _T_555; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_564 = $signed(spriteYRegs_38) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_565 = $signed(spriteYRegs_14) < $signed(_T_564); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_566 = _T_556 & $signed(spriteXRegs_38) < $signed(_T_99) & _T_565; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_571 = _T_566 & $signed(spriteYRegs_38) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire [10:0] _T_574 = $signed(spriteXRegs_39) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_575 = $signed(spriteXRegs_14) < $signed(_T_574); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_576 = spriteVisibleRegs_39 & _T_575; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_584 = $signed(spriteYRegs_39) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_585 = $signed(spriteYRegs_14) < $signed(_T_584); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_586 = _T_576 & $signed(spriteXRegs_39) < $signed(_T_99) & _T_585; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_591 = _T_586 & $signed(spriteYRegs_39) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire [10:0] _T_594 = $signed(spriteXRegs_40) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_595 = $signed(spriteXRegs_14) < $signed(_T_594); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_596 = spriteVisibleRegs_40 & _T_595; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_604 = $signed(spriteYRegs_40) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_605 = $signed(spriteYRegs_14) < $signed(_T_604); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_606 = _T_596 & $signed(spriteXRegs_40) < $signed(_T_99) & _T_605; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_611 = _T_606 & $signed(spriteYRegs_40) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire [10:0] _T_614 = $signed(spriteXRegs_41) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_615 = $signed(spriteXRegs_14) < $signed(_T_614); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_616 = spriteVisibleRegs_41 & _T_615; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_624 = $signed(spriteYRegs_41) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_625 = $signed(spriteYRegs_14) < $signed(_T_624); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_626 = _T_616 & $signed(spriteXRegs_41) < $signed(_T_99) & _T_625; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_631 = _T_626 & $signed(spriteYRegs_41) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire [10:0] _T_634 = $signed(spriteXRegs_42) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_635 = $signed(spriteXRegs_14) < $signed(_T_634); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_636 = spriteVisibleRegs_42 & _T_635; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_644 = $signed(spriteYRegs_42) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_645 = $signed(spriteYRegs_14) < $signed(_T_644); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_646 = _T_636 & $signed(spriteXRegs_42) < $signed(_T_99) & _T_645; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_651 = _T_646 & $signed(spriteYRegs_42) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire [10:0] _T_654 = $signed(spriteXRegs_43) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_655 = $signed(spriteXRegs_14) < $signed(_T_654); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_656 = spriteVisibleRegs_43 & _T_655; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_664 = $signed(spriteYRegs_43) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_665 = $signed(spriteYRegs_14) < $signed(_T_664); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_666 = _T_656 & $signed(spriteXRegs_43) < $signed(_T_99) & _T_665; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_671 = _T_666 & $signed(spriteYRegs_43) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire [10:0] _T_674 = $signed(spriteXRegs_44) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_675 = $signed(spriteXRegs_14) < $signed(_T_674); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_676 = spriteVisibleRegs_44 & _T_675; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_684 = $signed(spriteYRegs_44) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_685 = $signed(spriteYRegs_14) < $signed(_T_684); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_686 = _T_676 & $signed(spriteXRegs_44) < $signed(_T_99) & _T_685; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_691 = _T_686 & $signed(spriteYRegs_44) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire [10:0] _T_694 = $signed(spriteXRegs_45) + 11'sh20; // @[\\src\\main\\scala\\GameLogic.scala 445:49]
  wire  _T_695 = $signed(spriteXRegs_14) < $signed(_T_694); // @[\\src\\main\\scala\\GameLogic.scala 445:32]
  wire  _T_696 = spriteVisibleRegs_45 & _T_695; // @[\\src\\main\\scala\\GameLogic.scala 444:34]
  wire [9:0] _T_704 = $signed(spriteYRegs_45) + 10'shf; // @[\\src\\main\\scala\\GameLogic.scala 446:49]
  wire  _T_705 = $signed(spriteYRegs_14) < $signed(_T_704); // @[\\src\\main\\scala\\GameLogic.scala 446:32]
  wire  _T_706 = _T_696 & $signed(spriteXRegs_45) < $signed(_T_99) & _T_705; // @[\\src\\main\\scala\\GameLogic.scala 445:101]
  wire  _T_711 = _T_706 & $signed(spriteYRegs_45) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 446:57]
  wire  _GEN_1039 = _T_711 | (_T_691 | (_T_671 | (_T_651 | (_T_631 | (_T_611 | (_T_591 | (_T_571 | (_T_551 | (_T_531 |
    _GEN_1029))))))))); // @[\\src\\main\\scala\\GameLogic.scala 447:13 448:31]
  wire  _GEN_1040 = _T_89 ? _GEN_1039 : _GEN_1029; // @[\\src\\main\\scala\\GameLogic.scala 441:25]
  wire [10:0] _T_714 = $signed(spriteXRegs_13) + 11'sh16; // @[\\src\\main\\scala\\GameLogic.scala 456:44]
  wire  _T_715 = $signed(spriteXRegs_14) < $signed(_T_714); // @[\\src\\main\\scala\\GameLogic.scala 456:26]
  wire  _T_716 = spriteVisibleRegs_13 & _T_715; // @[\\src\\main\\scala\\GameLogic.scala 455:31]
  wire [9:0] _T_724 = $signed(spriteYRegs_13) + 10'sh16; // @[\\src\\main\\scala\\GameLogic.scala 457:44]
  wire  _T_725 = $signed(spriteYRegs_14) < $signed(_T_724); // @[\\src\\main\\scala\\GameLogic.scala 457:26]
  wire  _T_726 = _T_716 & $signed(spriteXRegs_13) < $signed(_T_99) & _T_725; // @[\\src\\main\\scala\\GameLogic.scala 456:97]
  wire  _T_731 = _T_726 & $signed(spriteYRegs_13) < $signed(_T_109); // @[\\src\\main\\scala\\GameLogic.scala 457:52]
  wire [2:0] _livesReg_T_1 = livesReg + 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 461:32]
  wire [2:0] _GEN_1041 = livesReg < 3'h3 ? _livesReg_T_1 : livesReg; // @[\\src\\main\\scala\\GameLogic.scala 460:30 461:20 223:25]
  wire [2:0] _GEN_1043 = _T_731 ? _GEN_1041 : livesReg; // @[\\src\\main\\scala\\GameLogic.scala 223:25 458:9]
  wire  _GEN_1044 = collisionDetected & _T_89 | isBlinking; // @[\\src\\main\\scala\\GameLogic.scala 466:46 467:20 242:27]
  wire [7:0] _GEN_1045 = collisionDetected & _T_89 ? 8'h0 : blinkCounter; // @[\\src\\main\\scala\\GameLogic.scala 466:46 468:22 240:29]
  wire [1:0] _GEN_1046 = collisionDetected & _T_89 ? 2'h0 : blinkTimes; // @[\\src\\main\\scala\\GameLogic.scala 466:46 469:20 241:27]
  wire  _GEN_1047 = blinkCounter < 8'h14 | _GEN_956; // @[\\src\\main\\scala\\GameLogic.scala 477:41 478:33]
  wire  _GEN_1048 = blinkCounter < 8'ha ? 1'h0 : _GEN_1047; // @[\\src\\main\\scala\\GameLogic.scala 475:35 476:33]
  wire [7:0] _blinkCounter_T_1 = blinkCounter + 8'h1; // @[\\src\\main\\scala\\GameLogic.scala 480:38]
  wire [1:0] _blinkTimes_T_1 = blinkTimes + 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 483:36]
  wire [7:0] _GEN_1049 = blinkCounter == 8'h14 ? 8'h0 : _blinkCounter_T_1; // @[\\src\\main\\scala\\GameLogic.scala 480:22 481:37 482:24]
  wire [1:0] _GEN_1050 = blinkCounter == 8'h14 ? _blinkTimes_T_1 : _GEN_1046; // @[\\src\\main\\scala\\GameLogic.scala 481:37 483:22]
  wire [2:0] _livesReg_T_3 = livesReg - 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 492:34]
  wire [2:0] _GEN_1051 = livesReg <= 3'h1 ? 3'h0 : _livesReg_T_3; // @[\\src\\main\\scala\\GameLogic.scala 488:33 489:22 492:22]
  wire [2:0] _GEN_1052 = livesReg <= 3'h1 ? 3'h6 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 488:33 490:22 113:25]
  wire  _GEN_1053 = blinkTimes == 2'h3 ? 1'h0 : _GEN_1044; // @[\\src\\main\\scala\\GameLogic.scala 485:34 486:22]
  wire  _GEN_1054 = blinkTimes == 2'h3 | _GEN_1048; // @[\\src\\main\\scala\\GameLogic.scala 485:34 487:33]
  wire [2:0] _GEN_1055 = blinkTimes == 2'h3 ? _GEN_1051 : _GEN_1043; // @[\\src\\main\\scala\\GameLogic.scala 485:34]
  wire [2:0] _GEN_1056 = blinkTimes == 2'h3 ? _GEN_1052 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 113:25 485:34]
  wire  _GEN_1057 = blinkTimes == 2'h3 ? 1'h0 : _GEN_1040; // @[\\src\\main\\scala\\GameLogic.scala 485:34 494:29]
  wire [2:0] _GEN_1063 = isBlinking ? _GEN_1056 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 473:24 113:25]
  reg [10:0] spriteXRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 513:35]
  reg [9:0] spriteYRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 514:35]
  reg [10:0] spriteXRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 515:35]
  reg [9:0] spriteYRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 516:35]
  reg [10:0] spriteXRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 517:35]
  reg [9:0] spriteYRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 518:35]
  wire [9:0] _starCnt_T_1 = starCnt + 10'h1; // @[\\src\\main\\scala\\GameLogic.scala 525:28]
  wire [10:0] _spriteXRegs_58_T_5 = $signed(spriteXRegs_58) + 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 533:44]
  wire [10:0] _spriteXRegs_59_T_5 = $signed(spriteXRegs_59) + 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 534:44]
  wire [10:0] _spriteXRegs_60_T_5 = $signed(spriteXRegs_60) + 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 535:44]
  wire [9:0] _spriteYRegs_58_T_5 = $signed(spriteYRegs_58) + 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 536:44]
  wire [9:0] _spriteYRegs_59_T_5 = $signed(spriteYRegs_59) + 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 537:44]
  wire [9:0] _spriteYRegs_60_T_5 = $signed(spriteYRegs_60) + 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 538:44]
  reg [10:0] spriteXRegs_58_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 541:35]
  reg [9:0] spriteYRegs_58_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 542:35]
  reg [10:0] spriteXRegs_59_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 543:35]
  reg [9:0] spriteYRegs_59_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 544:35]
  reg [10:0] spriteXRegs_60_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 545:35]
  reg [9:0] spriteYRegs_60_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 546:35]
  reg [10:0] spriteXRegs_58_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 569:35]
  reg [9:0] spriteYRegs_58_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 570:35]
  reg [10:0] spriteXRegs_59_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 571:35]
  reg [9:0] spriteYRegs_59_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 572:35]
  reg [10:0] spriteXRegs_60_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 573:35]
  reg [9:0] spriteYRegs_60_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 574:35]
  wire [9:0] _GEN_1066 = starCnt == 10'h168 ? 10'h0 : _starCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 596:37 597:17 599:17]
  wire  _GEN_1067 = starCnt == 10'h12c ? 1'h0 : sprite58ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 582:37 583:35 169:42]
  wire  _GEN_1068 = starCnt == 10'h12c ? 1'h0 : sprite59ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 582:37 584:35 171:42]
  wire  _GEN_1069 = starCnt == 10'h12c ? 1'h0 : sprite60ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 582:37 585:35 173:42]
  wire  _GEN_1070 = starCnt == 10'h12c ? 1'h0 : sprite58ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 582:37 586:33 170:40]
  wire  _GEN_1071 = starCnt == 10'h12c ? 1'h0 : sprite59ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 582:37 587:33 172:40]
  wire  _GEN_1072 = starCnt == 10'h12c ? 1'h0 : sprite60ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 582:37 588:33 174:40]
  wire [10:0] _GEN_1073 = starCnt == 10'h12c ? $signed(_spriteXRegs_58_T_5) : $signed(_GEN_102); // @[\\src\\main\\scala\\GameLogic.scala 582:37 589:25]
  wire [10:0] _GEN_1074 = starCnt == 10'h12c ? $signed(_spriteXRegs_59_T_5) : $signed(_GEN_104); // @[\\src\\main\\scala\\GameLogic.scala 582:37 590:25]
  wire [10:0] _GEN_1075 = starCnt == 10'h12c ? $signed(_spriteXRegs_60_T_5) : $signed(_GEN_106); // @[\\src\\main\\scala\\GameLogic.scala 582:37 591:25]
  wire [9:0] _GEN_1076 = starCnt == 10'h12c ? $signed(_spriteYRegs_58_T_5) : $signed(_GEN_103); // @[\\src\\main\\scala\\GameLogic.scala 582:37 592:25]
  wire [9:0] _GEN_1077 = starCnt == 10'h12c ? $signed(_spriteYRegs_59_T_5) : $signed(_GEN_105); // @[\\src\\main\\scala\\GameLogic.scala 582:37 593:25]
  wire [9:0] _GEN_1078 = starCnt == 10'h12c ? $signed(_spriteYRegs_60_T_5) : $signed(_GEN_107); // @[\\src\\main\\scala\\GameLogic.scala 582:37 594:25]
  wire [9:0] _GEN_1079 = starCnt == 10'h12c ? _starCnt_T_1 : _GEN_1066; // @[\\src\\main\\scala\\GameLogic.scala 582:37 595:17]
  wire [10:0] _GEN_1080 = starCnt == 10'hf0 ? $signed(spriteXRegs_58_REG_2) : $signed(_GEN_1073); // @[\\src\\main\\scala\\GameLogic.scala 568:37 569:25]
  wire [9:0] _GEN_1081 = starCnt == 10'hf0 ? $signed(spriteYRegs_58_REG_2) : $signed(_GEN_1076); // @[\\src\\main\\scala\\GameLogic.scala 568:37 570:25]
  wire [10:0] _GEN_1082 = starCnt == 10'hf0 ? $signed(spriteXRegs_59_REG_2) : $signed(_GEN_1074); // @[\\src\\main\\scala\\GameLogic.scala 568:37 571:25]
  wire [9:0] _GEN_1083 = starCnt == 10'hf0 ? $signed(spriteYRegs_59_REG_2) : $signed(_GEN_1077); // @[\\src\\main\\scala\\GameLogic.scala 568:37 572:25]
  wire [10:0] _GEN_1084 = starCnt == 10'hf0 ? $signed(spriteXRegs_60_REG_2) : $signed(_GEN_1075); // @[\\src\\main\\scala\\GameLogic.scala 568:37 573:25]
  wire [9:0] _GEN_1085 = starCnt == 10'hf0 ? $signed(spriteYRegs_60_REG_2) : $signed(_GEN_1078); // @[\\src\\main\\scala\\GameLogic.scala 568:37 574:25]
  wire  _GEN_1086 = starCnt == 10'hf0 | _GEN_1067; // @[\\src\\main\\scala\\GameLogic.scala 568:37 575:35]
  wire  _GEN_1087 = starCnt == 10'hf0 | _GEN_1068; // @[\\src\\main\\scala\\GameLogic.scala 568:37 576:35]
  wire  _GEN_1088 = starCnt == 10'hf0 | _GEN_1069; // @[\\src\\main\\scala\\GameLogic.scala 568:37 577:35]
  wire  _GEN_1089 = starCnt == 10'hf0 | _GEN_1070; // @[\\src\\main\\scala\\GameLogic.scala 568:37 578:33]
  wire  _GEN_1090 = starCnt == 10'hf0 | _GEN_1071; // @[\\src\\main\\scala\\GameLogic.scala 568:37 579:33]
  wire  _GEN_1091 = starCnt == 10'hf0 | _GEN_1072; // @[\\src\\main\\scala\\GameLogic.scala 568:37 580:33]
  wire [9:0] _GEN_1092 = starCnt == 10'hf0 ? _starCnt_T_1 : _GEN_1079; // @[\\src\\main\\scala\\GameLogic.scala 568:37 581:17]
  wire  _GEN_1093 = starCnt == 10'hb4 ? 1'h0 : _GEN_1086; // @[\\src\\main\\scala\\GameLogic.scala 554:37 555:35]
  wire  _GEN_1094 = starCnt == 10'hb4 ? 1'h0 : _GEN_1087; // @[\\src\\main\\scala\\GameLogic.scala 554:37 556:35]
  wire  _GEN_1095 = starCnt == 10'hb4 ? 1'h0 : _GEN_1088; // @[\\src\\main\\scala\\GameLogic.scala 554:37 557:35]
  wire  _GEN_1096 = starCnt == 10'hb4 ? 1'h0 : _GEN_1089; // @[\\src\\main\\scala\\GameLogic.scala 554:37 558:33]
  wire  _GEN_1097 = starCnt == 10'hb4 ? 1'h0 : _GEN_1090; // @[\\src\\main\\scala\\GameLogic.scala 554:37 559:33]
  wire  _GEN_1098 = starCnt == 10'hb4 ? 1'h0 : _GEN_1091; // @[\\src\\main\\scala\\GameLogic.scala 554:37 560:33]
  wire [10:0] _GEN_1099 = starCnt == 10'hb4 ? $signed(_spriteXRegs_58_T_5) : $signed(_GEN_1080); // @[\\src\\main\\scala\\GameLogic.scala 554:37 561:25]
  wire [10:0] _GEN_1100 = starCnt == 10'hb4 ? $signed(_spriteXRegs_59_T_5) : $signed(_GEN_1082); // @[\\src\\main\\scala\\GameLogic.scala 554:37 562:25]
  wire [10:0] _GEN_1101 = starCnt == 10'hb4 ? $signed(_spriteXRegs_60_T_5) : $signed(_GEN_1084); // @[\\src\\main\\scala\\GameLogic.scala 554:37 563:25]
  wire [9:0] _GEN_1102 = starCnt == 10'hb4 ? $signed(_spriteYRegs_58_T_5) : $signed(_GEN_1081); // @[\\src\\main\\scala\\GameLogic.scala 554:37 564:25]
  wire [9:0] _GEN_1103 = starCnt == 10'hb4 ? $signed(_spriteYRegs_59_T_5) : $signed(_GEN_1083); // @[\\src\\main\\scala\\GameLogic.scala 554:37 565:25]
  wire [9:0] _GEN_1104 = starCnt == 10'hb4 ? $signed(_spriteYRegs_60_T_5) : $signed(_GEN_1085); // @[\\src\\main\\scala\\GameLogic.scala 554:37 566:25]
  wire [9:0] _GEN_1105 = starCnt == 10'hb4 ? _starCnt_T_1 : _GEN_1092; // @[\\src\\main\\scala\\GameLogic.scala 554:37 567:17]
  wire [10:0] _GEN_1106 = starCnt == 10'h78 ? $signed(spriteXRegs_58_REG_1) : $signed(_GEN_1099); // @[\\src\\main\\scala\\GameLogic.scala 540:37 541:25]
  wire [9:0] _GEN_1107 = starCnt == 10'h78 ? $signed(spriteYRegs_58_REG_1) : $signed(_GEN_1102); // @[\\src\\main\\scala\\GameLogic.scala 540:37 542:25]
  wire [10:0] _GEN_1108 = starCnt == 10'h78 ? $signed(spriteXRegs_59_REG_1) : $signed(_GEN_1100); // @[\\src\\main\\scala\\GameLogic.scala 540:37 543:25]
  wire [9:0] _GEN_1109 = starCnt == 10'h78 ? $signed(spriteYRegs_59_REG_1) : $signed(_GEN_1103); // @[\\src\\main\\scala\\GameLogic.scala 540:37 544:25]
  wire [10:0] _GEN_1110 = starCnt == 10'h78 ? $signed(spriteXRegs_60_REG_1) : $signed(_GEN_1101); // @[\\src\\main\\scala\\GameLogic.scala 540:37 545:25]
  wire [9:0] _GEN_1111 = starCnt == 10'h78 ? $signed(spriteYRegs_60_REG_1) : $signed(_GEN_1104); // @[\\src\\main\\scala\\GameLogic.scala 540:37 546:25]
  wire  _GEN_1112 = starCnt == 10'h78 | _GEN_1093; // @[\\src\\main\\scala\\GameLogic.scala 540:37 547:35]
  wire  _GEN_1113 = starCnt == 10'h78 | _GEN_1094; // @[\\src\\main\\scala\\GameLogic.scala 540:37 548:35]
  wire  _GEN_1114 = starCnt == 10'h78 | _GEN_1095; // @[\\src\\main\\scala\\GameLogic.scala 540:37 549:35]
  wire  _GEN_1115 = starCnt == 10'h78 | _GEN_1096; // @[\\src\\main\\scala\\GameLogic.scala 540:37 550:33]
  wire  _GEN_1116 = starCnt == 10'h78 | _GEN_1097; // @[\\src\\main\\scala\\GameLogic.scala 540:37 551:33]
  wire  _GEN_1117 = starCnt == 10'h78 | _GEN_1098; // @[\\src\\main\\scala\\GameLogic.scala 540:37 552:33]
  wire [9:0] _GEN_1118 = starCnt == 10'h78 ? _starCnt_T_1 : _GEN_1105; // @[\\src\\main\\scala\\GameLogic.scala 540:37 553:17]
  wire  _GEN_1119 = starCnt == 10'h3c ? 1'h0 : _GEN_1112; // @[\\src\\main\\scala\\GameLogic.scala 526:36 527:35]
  wire  _GEN_1120 = starCnt == 10'h3c ? 1'h0 : _GEN_1113; // @[\\src\\main\\scala\\GameLogic.scala 526:36 528:35]
  wire  _GEN_1121 = starCnt == 10'h3c ? 1'h0 : _GEN_1114; // @[\\src\\main\\scala\\GameLogic.scala 526:36 529:35]
  wire  _GEN_1122 = starCnt == 10'h3c ? 1'h0 : _GEN_1115; // @[\\src\\main\\scala\\GameLogic.scala 526:36 530:33]
  wire  _GEN_1123 = starCnt == 10'h3c ? 1'h0 : _GEN_1116; // @[\\src\\main\\scala\\GameLogic.scala 526:36 531:33]
  wire  _GEN_1124 = starCnt == 10'h3c ? 1'h0 : _GEN_1117; // @[\\src\\main\\scala\\GameLogic.scala 526:36 532:33]
  wire [10:0] _GEN_1125 = starCnt == 10'h3c ? $signed(_spriteXRegs_58_T_5) : $signed(_GEN_1106); // @[\\src\\main\\scala\\GameLogic.scala 526:36 533:25]
  wire [10:0] _GEN_1126 = starCnt == 10'h3c ? $signed(_spriteXRegs_59_T_5) : $signed(_GEN_1108); // @[\\src\\main\\scala\\GameLogic.scala 526:36 534:25]
  wire [10:0] _GEN_1127 = starCnt == 10'h3c ? $signed(_spriteXRegs_60_T_5) : $signed(_GEN_1110); // @[\\src\\main\\scala\\GameLogic.scala 526:36 535:25]
  wire [9:0] _GEN_1128 = starCnt == 10'h3c ? $signed(_spriteYRegs_58_T_5) : $signed(_GEN_1107); // @[\\src\\main\\scala\\GameLogic.scala 526:36 536:25]
  wire [9:0] _GEN_1129 = starCnt == 10'h3c ? $signed(_spriteYRegs_59_T_5) : $signed(_GEN_1109); // @[\\src\\main\\scala\\GameLogic.scala 526:36 537:25]
  wire [9:0] _GEN_1130 = starCnt == 10'h3c ? $signed(_spriteYRegs_60_T_5) : $signed(_GEN_1111); // @[\\src\\main\\scala\\GameLogic.scala 526:36 538:25]
  wire [9:0] _GEN_1131 = starCnt == 10'h3c ? _starCnt_T_1 : _GEN_1118; // @[\\src\\main\\scala\\GameLogic.scala 526:36 539:17]
  wire  _GEN_1138 = starCnt == 10'h0 | _GEN_1119; // @[\\src\\main\\scala\\GameLogic.scala 512:29 519:35]
  wire  _GEN_1139 = starCnt == 10'h0 | _GEN_1120; // @[\\src\\main\\scala\\GameLogic.scala 512:29 520:35]
  wire  _GEN_1140 = starCnt == 10'h0 | _GEN_1121; // @[\\src\\main\\scala\\GameLogic.scala 512:29 521:35]
  wire  _GEN_1141 = starCnt == 10'h0 | _GEN_1122; // @[\\src\\main\\scala\\GameLogic.scala 512:29 522:33]
  wire  _GEN_1142 = starCnt == 10'h0 | _GEN_1123; // @[\\src\\main\\scala\\GameLogic.scala 512:29 523:33]
  wire  _GEN_1143 = starCnt == 10'h0 | _GEN_1124; // @[\\src\\main\\scala\\GameLogic.scala 512:29 524:33]
  wire  _T_754 = $signed(spriteYRegs_3) > 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 620:81]
  wire  _T_756 = $signed(spriteYRegs_3) < 10'sh14c; // @[\\src\\main\\scala\\GameLogic.scala 620:107]
  wire  _T_757 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c; // @[\\src\\main\\scala\\GameLogic.scala 620:89]
  wire [1:0] _GEN_1146 = io_btnC ? 2'h1 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 623:25 624:20 212:23]
  wire [2:0] _GEN_1147 = io_btnC ? 3'h3 : 3'h4; // @[\\src\\main\\scala\\GameLogic.scala 623:25 625:22 627:22]
  wire  _T_764 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_754 & _T_756; // @[\\src\\main\\scala\\GameLogic.scala 629:95]
  wire [1:0] _GEN_1148 = io_btnC ? 2'h2 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 632:25 633:20 212:23]
  wire  _T_771 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_754 & _T_756; // @[\\src\\main\\scala\\GameLogic.scala 638:95]
  wire [1:0] _GEN_1149 = io_btnC ? 2'h3 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 641:25 642:20 212:23]
  wire  _GEN_1150 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_754 & _T_756 ? 1'h0 : 1'h1
    ; // @[\\src\\main\\scala\\GameLogic.scala 638:122 617:31 639:33]
  wire [1:0] _GEN_1152 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_754 & _T_756 ?
    _GEN_1149 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 638:122 212:23]
  wire [2:0] _GEN_1153 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_754 & _T_756 ?
    _GEN_1147 : 3'h4; // @[\\src\\main\\scala\\GameLogic.scala 638:122 648:20]
  wire  _GEN_1154 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_754 & _T_756 ? 1'h0 : 1'h1
    ; // @[\\src\\main\\scala\\GameLogic.scala 629:122 615:30 630:32]
  wire [1:0] _GEN_1156 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_754 & _T_756 ?
    _GEN_1148 : _GEN_1152; // @[\\src\\main\\scala\\GameLogic.scala 629:122]
  wire [2:0] _GEN_1157 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_754 & _T_756 ?
    _GEN_1147 : _GEN_1153; // @[\\src\\main\\scala\\GameLogic.scala 629:122]
  wire  _GEN_1158 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_754 & _T_756 | _GEN_1150; // @[\\src\\main\\scala\\GameLogic.scala 629:122 617:31]
  wire  _GEN_1159 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_754 & _T_756 ? 1'h0 :
    _T_771; // @[\\src\\main\\scala\\GameLogic.scala 629:122 618:31]
  wire  _GEN_1160 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 620:116 613:30 621:32]
  wire [1:0] _GEN_1162 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3)
     > 10'sh12c & $signed(spriteYRegs_3) < 10'sh14c ? _GEN_1146 : _GEN_1156; // @[\\src\\main\\scala\\GameLogic.scala 620:116]
  wire [2:0] _GEN_1163 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3)
     > 10'sh12c & $signed(spriteYRegs_3) < 10'sh14c ? _GEN_1147 : _GEN_1157; // @[\\src\\main\\scala\\GameLogic.scala 620:116]
  wire  _GEN_1164 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c | _GEN_1154; // @[\\src\\main\\scala\\GameLogic.scala 620:116 615:30]
  wire  _GEN_1165 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c ? 1'h0 : _T_764; // @[\\src\\main\\scala\\GameLogic.scala 620:116 616:31]
  wire  _GEN_1166 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c | _GEN_1158; // @[\\src\\main\\scala\\GameLogic.scala 620:116 617:31]
  wire  _GEN_1167 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c ? 1'h0 : _GEN_1159; // @[\\src\\main\\scala\\GameLogic.scala 620:116 618:31]
  wire [2:0] _GEN_1168 = _T ? 3'h4 : _GEN_1163; // @[\\src\\main\\scala\\GameLogic.scala 608:28 609:18]
  wire  _GEN_1169 = _T ? spriteVisibleRegs_3 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 608:28 125:34 612:30]
  wire  _GEN_1170 = _T ? spriteVisibleRegs_7 : _GEN_1160; // @[\\src\\main\\scala\\GameLogic.scala 608:28 125:34]
  wire  _GEN_1171 = _T ? spriteVisibleRegs_8 : _T_757; // @[\\src\\main\\scala\\GameLogic.scala 608:28 125:34]
  wire  _GEN_1172 = _T ? spriteVisibleRegs_9 : _GEN_1164; // @[\\src\\main\\scala\\GameLogic.scala 608:28 125:34]
  wire  _GEN_1173 = _T ? spriteVisibleRegs_10 : _GEN_1165; // @[\\src\\main\\scala\\GameLogic.scala 608:28 125:34]
  wire  _GEN_1174 = _T ? spriteVisibleRegs_11 : _GEN_1166; // @[\\src\\main\\scala\\GameLogic.scala 608:28 125:34]
  wire  _GEN_1175 = _T ? spriteVisibleRegs_12 : _GEN_1167; // @[\\src\\main\\scala\\GameLogic.scala 608:28 125:34]
  wire [1:0] _GEN_1176 = _T ? lvlReg : _GEN_1162; // @[\\src\\main\\scala\\GameLogic.scala 212:23 608:28]
  wire [9:0] _GEN_1177 = _T_82 ? 10'h280 : viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 676:34 677:21 202:28]
  wire [8:0] _GEN_1178 = _T_82 ? 9'h1e0 : viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 676:34 678:21 203:28]
  wire [9:0] _GEN_1179 = _T_75 ? 10'h0 : _GEN_1177; // @[\\src\\main\\scala\\GameLogic.scala 673:34 674:21]
  wire [8:0] _GEN_1180 = _T_75 ? 9'h1e0 : _GEN_1178; // @[\\src\\main\\scala\\GameLogic.scala 673:34 675:21]
  wire [9:0] _GEN_1181 = _T_68 ? 10'h280 : _GEN_1179; // @[\\src\\main\\scala\\GameLogic.scala 670:28 671:21]
  wire [8:0] _GEN_1182 = _T_68 ? 9'h0 : _GEN_1180; // @[\\src\\main\\scala\\GameLogic.scala 670:28 672:21]
  wire [9:0] _spriteYRegs_14_T_2 = $signed(spriteYRegs_14) + 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 688:48]
  wire [9:0] _GEN_1183 = $signed(spriteYRegs_14) < 10'sh1c0 ? $signed(_spriteYRegs_14_T_2) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 687:48 688:29]
  wire [9:0] _spriteYRegs_14_T_5 = $signed(spriteYRegs_14) - 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 692:48]
  wire [9:0] _GEN_1184 = $signed(spriteYRegs_14) > 10'sh20 ? $signed(_spriteYRegs_14_T_5) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 691:40 692:29]
  wire [9:0] _GEN_1185 = io_btnU ? $signed(_GEN_1184) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 690:29]
  wire [9:0] _GEN_1186 = io_btnD ? $signed(_GEN_1183) : $signed(_GEN_1185); // @[\\src\\main\\scala\\GameLogic.scala 686:22]
  wire [9:0] _spriteYRegs_3_T_2 = $signed(spriteYRegs_3) + 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 699:46]
  wire [9:0] _GEN_1187 = $signed(spriteYRegs_3) < 10'sh1c0 ? $signed(_spriteYRegs_3_T_2) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 698:47 699:28]
  wire [9:0] _spriteYRegs_3_T_5 = $signed(spriteYRegs_3) - 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 703:46]
  wire [9:0] _GEN_1188 = $signed(spriteYRegs_3) > 10'sh20 ? $signed(_spriteYRegs_3_T_5) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 702:39 703:28]
  wire [9:0] _GEN_1189 = io_btnU ? $signed(_GEN_1188) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 701:29]
  wire [9:0] _GEN_1190 = io_btnD ? $signed(_GEN_1187) : $signed(_GEN_1189); // @[\\src\\main\\scala\\GameLogic.scala 697:22]
  wire [10:0] _spriteXRegs_3_T_2 = $signed(spriteXRegs_3) + 11'sh2; // @[\\src\\main\\scala\\GameLogic.scala 708:46]
  wire [10:0] _GEN_1191 = $signed(spriteXRegs_3) < 11'sh260 ? $signed(_spriteXRegs_3_T_2) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 707:47 708:28]
  wire [10:0] _spriteXRegs_3_T_5 = $signed(spriteXRegs_3) - 11'sh2; // @[\\src\\main\\scala\\GameLogic.scala 712:46]
  wire [10:0] _GEN_1192 = $signed(spriteXRegs_3) > 11'sh20 ? $signed(_spriteXRegs_3_T_5) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 711:39 712:28]
  wire [10:0] _GEN_1193 = io_btnL ? $signed(_GEN_1192) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 710:29]
  wire [10:0] _GEN_1194 = io_btnR ? $signed(_GEN_1191) : $signed(_GEN_1193); // @[\\src\\main\\scala\\GameLogic.scala 706:23]
  wire [9:0] _GEN_1195 = _T ? $signed(_GEN_1186) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 685:28]
  wire [9:0] _GEN_1196 = _T ? $signed(_GEN_1) : $signed(_GEN_1190); // @[\\src\\main\\scala\\GameLogic.scala 685:28]
  wire [10:0] _GEN_1197 = _T ? $signed(_GEN_0) : $signed(_GEN_1194); // @[\\src\\main\\scala\\GameLogic.scala 685:28]
  wire [2:0] _GEN_1198 = $signed(spriteXRegs_3) > 11'sh104 & $signed(spriteXRegs_3) < 11'sh17c & $signed(spriteYRegs_3)
     > 10'sh122 & $signed(spriteYRegs_3) < 10'sh154 & io_btnC ? 3'h2 : 3'h4; // @[\\src\\main\\scala\\GameLogic.scala 741:125 742:18 747:18]
  wire [1:0] _GEN_1199 = $signed(spriteXRegs_3) > 11'sh104 & $signed(spriteXRegs_3) < 11'sh17c & $signed(spriteYRegs_3)
     > 10'sh122 & $signed(spriteYRegs_3) < 10'sh154 & io_btnC ? 2'h0 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 741:125 743:16 212:23]
  wire [2:0] _GEN_1200 = $signed(spriteXRegs_3) > 11'sh104 & $signed(spriteXRegs_3) < 11'sh17c & $signed(spriteYRegs_3)
     > 10'sh122 & $signed(spriteYRegs_3) < 10'sh154 & io_btnC ? 3'h3 : livesReg; // @[\\src\\main\\scala\\GameLogic.scala 741:125 744:18 223:25]
  wire [2:0] _GEN_1203 = 3'h5 == stateReg ? 3'h0 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 279:20 752:16 113:25]
  wire  _GEN_1204 = 3'h6 == stateReg ? 1'h0 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 279:20 720:29 125:34]
  wire  _GEN_1205 = 3'h6 == stateReg | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 279:20 723:29 125:34]
  wire  _GEN_1206 = 3'h6 == stateReg | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 279:20 724:29 125:34]
  wire  _GEN_1207 = 3'h6 == stateReg | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 279:20 725:29 125:34]
  wire  _GEN_1208 = 3'h6 == stateReg | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 279:20 726:29 125:34]
  wire  _GEN_1209 = 3'h6 == stateReg | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 279:20 727:29 125:34]
  wire  _GEN_1210 = 3'h6 == stateReg | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 279:20 728:29 125:34]
  wire  _GEN_1211 = 3'h6 == stateReg | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 279:20 730:29 125:34]
  wire  _GEN_1212 = 3'h6 == stateReg | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 279:20 731:29 125:34]
  wire  _GEN_1213 = 3'h6 == stateReg | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 279:20 732:29 125:34]
  wire  _GEN_1214 = 3'h6 == stateReg | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 279:20 733:29 125:34]
  wire  _GEN_1215 = 3'h6 == stateReg | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 279:20 734:29 125:34]
  wire  _GEN_1216 = 3'h6 == stateReg | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 279:20 735:29 125:34]
  wire  _GEN_1217 = 3'h6 == stateReg | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 279:20 738:29 125:34]
  wire [2:0] _GEN_1218 = 3'h6 == stateReg ? _GEN_1198 : _GEN_1203; // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [1:0] _GEN_1219 = 3'h6 == stateReg ? _GEN_1199 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 279:20 212:23]
  wire [2:0] _GEN_1220 = 3'h6 == stateReg ? _GEN_1200 : livesReg; // @[\\src\\main\\scala\\GameLogic.scala 279:20 223:25]
  wire  _GEN_1222 = 3'h6 == stateReg ? 1'h0 : 3'h5 == stateReg; // @[\\src\\main\\scala\\GameLogic.scala 279:20 100:22]
  wire [9:0] _GEN_1223 = 3'h4 == stateReg ? $signed(_GEN_1195) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [9:0] _GEN_1224 = 3'h4 == stateReg ? $signed(_GEN_1196) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [10:0] _GEN_1225 = 3'h4 == stateReg ? $signed(_GEN_1197) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [2:0] _GEN_1226 = 3'h4 == stateReg ? 3'h5 : _GEN_1218; // @[\\src\\main\\scala\\GameLogic.scala 279:20 716:16]
  wire  _GEN_1227 = 3'h4 == stateReg ? spriteVisibleRegs_14 : _GEN_1204; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1228 = 3'h4 == stateReg ? spriteVisibleRegs_46 : _GEN_1205; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1229 = 3'h4 == stateReg ? spriteVisibleRegs_47 : _GEN_1206; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1230 = 3'h4 == stateReg ? spriteVisibleRegs_48 : _GEN_1207; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1231 = 3'h4 == stateReg ? spriteVisibleRegs_49 : _GEN_1208; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1232 = 3'h4 == stateReg ? spriteVisibleRegs_50 : _GEN_1209; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1233 = 3'h4 == stateReg ? spriteVisibleRegs_51 : _GEN_1210; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1234 = 3'h4 == stateReg ? spriteVisibleRegs_52 : _GEN_1211; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1235 = 3'h4 == stateReg ? spriteVisibleRegs_53 : _GEN_1212; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1236 = 3'h4 == stateReg ? spriteVisibleRegs_54 : _GEN_1213; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1237 = 3'h4 == stateReg ? spriteVisibleRegs_55 : _GEN_1214; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1238 = 3'h4 == stateReg ? spriteVisibleRegs_56 : _GEN_1215; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1239 = 3'h4 == stateReg ? spriteVisibleRegs_57 : _GEN_1216; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1240 = 3'h4 == stateReg ? spriteVisibleRegs_3 : _GEN_1217; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire [1:0] _GEN_1241 = 3'h4 == stateReg ? lvlReg : _GEN_1219; // @[\\src\\main\\scala\\GameLogic.scala 279:20 212:23]
  wire [2:0] _GEN_1242 = 3'h4 == stateReg ? livesReg : _GEN_1220; // @[\\src\\main\\scala\\GameLogic.scala 279:20 223:25]
  wire  _GEN_1244 = 3'h4 == stateReg ? 1'h0 : _GEN_1222; // @[\\src\\main\\scala\\GameLogic.scala 279:20 100:22]
  wire [5:0] _GEN_1245 = 3'h3 == stateReg ? 6'h0 : nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 279:20 654:25 233:34]
  wire [7:0] _GEN_1246 = 3'h3 == stateReg ? 8'h0 : spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 279:20 655:25 232:34]
  wire [10:0] _GEN_1247 = 3'h3 == stateReg ? $signed(11'sh260) : $signed(_GEN_16); // @[\\src\\main\\scala\\GameLogic.scala 279:20 657:23]
  wire [9:0] _GEN_1248 = 3'h3 == stateReg ? $signed(10'sh140) : $signed(_GEN_1223); // @[\\src\\main\\scala\\GameLogic.scala 279:20 658:23]
  wire  _GEN_1249 = 3'h3 == stateReg ? 1'h0 : _GEN_1240; // @[\\src\\main\\scala\\GameLogic.scala 279:20 659:28]
  wire  _GEN_1250 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 279:20 660:28 125:34]
  wire  _GEN_1251 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 279:20 661:28 125:34]
  wire  _GEN_1252 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 279:20 662:28 125:34]
  wire  _GEN_1253 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 279:20 663:29 125:34]
  wire  _GEN_1254 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 279:20 664:29 125:34]
  wire  _GEN_1255 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 279:20 665:29 125:34]
  wire  _GEN_1256 = 3'h3 == stateReg | _GEN_1227; // @[\\src\\main\\scala\\GameLogic.scala 279:20 666:29]
  wire  _GEN_1257 = 3'h3 == stateReg | _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 279:20 667:29]
  wire  _GEN_1258 = 3'h3 == stateReg | _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 279:20 668:29]
  wire  _GEN_1259 = 3'h3 == stateReg | _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 279:20 669:29]
  wire [9:0] _GEN_1260 = 3'h3 == stateReg ? _GEN_1181 : viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 279:20 202:28]
  wire [8:0] _GEN_1261 = 3'h3 == stateReg ? _GEN_1182 : viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 279:20 203:28]
  wire [2:0] _GEN_1262 = 3'h3 == stateReg ? 3'h4 : _GEN_1226; // @[\\src\\main\\scala\\GameLogic.scala 279:20 680:16]
  wire [9:0] _GEN_1263 = 3'h3 == stateReg ? $signed(_GEN_1) : $signed(_GEN_1224); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [10:0] _GEN_1264 = 3'h3 == stateReg ? $signed(_GEN_0) : $signed(_GEN_1225); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1265 = 3'h3 == stateReg ? spriteVisibleRegs_46 : _GEN_1228; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1266 = 3'h3 == stateReg ? spriteVisibleRegs_47 : _GEN_1229; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1267 = 3'h3 == stateReg ? spriteVisibleRegs_48 : _GEN_1230; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1268 = 3'h3 == stateReg ? spriteVisibleRegs_49 : _GEN_1231; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1269 = 3'h3 == stateReg ? spriteVisibleRegs_50 : _GEN_1232; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1270 = 3'h3 == stateReg ? spriteVisibleRegs_51 : _GEN_1233; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1271 = 3'h3 == stateReg ? spriteVisibleRegs_52 : _GEN_1234; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1272 = 3'h3 == stateReg ? spriteVisibleRegs_53 : _GEN_1235; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1273 = 3'h3 == stateReg ? spriteVisibleRegs_54 : _GEN_1236; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1274 = 3'h3 == stateReg ? spriteVisibleRegs_55 : _GEN_1237; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1275 = 3'h3 == stateReg ? spriteVisibleRegs_56 : _GEN_1238; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire  _GEN_1276 = 3'h3 == stateReg ? spriteVisibleRegs_57 : _GEN_1239; // @[\\src\\main\\scala\\GameLogic.scala 279:20 125:34]
  wire [1:0] _GEN_1277 = 3'h3 == stateReg ? lvlReg : _GEN_1241; // @[\\src\\main\\scala\\GameLogic.scala 279:20 212:23]
  wire [2:0] _GEN_1278 = 3'h3 == stateReg ? livesReg : _GEN_1242; // @[\\src\\main\\scala\\GameLogic.scala 279:20 223:25]
  wire  _GEN_1280 = 3'h3 == stateReg ? 1'h0 : _GEN_1244; // @[\\src\\main\\scala\\GameLogic.scala 279:20 100:22]
  wire  _GEN_1316 = 3'h2 == stateReg ? 1'h0 : _GEN_1280; // @[\\src\\main\\scala\\GameLogic.scala 279:20 100:22]
  wire [26:0] _GEN_1319 = 3'h1 == stateReg ? $signed(_GEN_283) : $signed({{16{_GEN_18[10]}},_GEN_18}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1322 = 3'h1 == stateReg ? _GEN_286 : spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1324 = 3'h1 == stateReg ? $signed(_GEN_288) : $signed({{16{_GEN_20[10]}},_GEN_20}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1327 = 3'h1 == stateReg ? _GEN_291 : spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1329 = 3'h1 == stateReg ? $signed(_GEN_293) : $signed({{16{_GEN_22[10]}},_GEN_22}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1332 = 3'h1 == stateReg ? _GEN_296 : spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1334 = 3'h1 == stateReg ? $signed(_GEN_298) : $signed({{16{_GEN_24[10]}},_GEN_24}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1337 = 3'h1 == stateReg ? _GEN_301 : spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1339 = 3'h1 == stateReg ? $signed(_GEN_303) : $signed({{16{_GEN_26[10]}},_GEN_26}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1342 = 3'h1 == stateReg ? _GEN_306 : spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1344 = 3'h1 == stateReg ? $signed(_GEN_308) : $signed({{16{_GEN_28[10]}},_GEN_28}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1347 = 3'h1 == stateReg ? _GEN_311 : spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1349 = 3'h1 == stateReg ? $signed(_GEN_313) : $signed({{16{_GEN_30[10]}},_GEN_30}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1352 = 3'h1 == stateReg ? _GEN_316 : spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1354 = 3'h1 == stateReg ? $signed(_GEN_318) : $signed({{16{_GEN_32[10]}},_GEN_32}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1357 = 3'h1 == stateReg ? _GEN_321 : spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1359 = 3'h1 == stateReg ? $signed(_GEN_323) : $signed({{16{_GEN_34[10]}},_GEN_34}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1362 = 3'h1 == stateReg ? _GEN_326 : spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1364 = 3'h1 == stateReg ? $signed(_GEN_328) : $signed({{16{_GEN_36[10]}},_GEN_36}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1367 = 3'h1 == stateReg ? _GEN_331 : spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  wire [26:0] _GEN_1369 = 3'h1 == stateReg ? $signed(_GEN_333) : $signed({{16{_GEN_38[10]}},_GEN_38}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1373 = 3'h1 == stateReg ? $signed(_GEN_337) : $signed({{16{_GEN_40[10]}},_GEN_40}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1377 = 3'h1 == stateReg ? $signed(_GEN_341) : $signed({{16{_GEN_42[10]}},_GEN_42}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1381 = 3'h1 == stateReg ? $signed(_GEN_345) : $signed({{16{_GEN_44[10]}},_GEN_44}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1385 = 3'h1 == stateReg ? $signed(_GEN_349) : $signed({{16{_GEN_46[10]}},_GEN_46}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1389 = 3'h1 == stateReg ? $signed(_GEN_353) : $signed({{16{_GEN_48[10]}},_GEN_48}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1393 = 3'h1 == stateReg ? $signed(_GEN_357) : $signed({{16{_GEN_50[10]}},_GEN_50}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1397 = 3'h1 == stateReg ? $signed(_GEN_361) : $signed({{16{_GEN_52[10]}},_GEN_52}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1401 = 3'h1 == stateReg ? $signed(_GEN_365) : $signed({{16{_GEN_54[10]}},_GEN_54}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1405 = 3'h1 == stateReg ? $signed(_GEN_369) : $signed({{16{_GEN_56[10]}},_GEN_56}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1409 = 3'h1 == stateReg ? $signed(_GEN_373) : $signed({{16{_GEN_58[10]}},_GEN_58}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1413 = 3'h1 == stateReg ? $signed(_GEN_377) : $signed({{16{_GEN_60[10]}},_GEN_60}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1417 = 3'h1 == stateReg ? $signed(_GEN_381) : $signed({{16{_GEN_62[10]}},_GEN_62}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1421 = 3'h1 == stateReg ? $signed(_GEN_385) : $signed({{16{_GEN_64[10]}},_GEN_64}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1425 = 3'h1 == stateReg ? $signed(_GEN_389) : $signed({{16{_GEN_66[10]}},_GEN_66}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1429 = 3'h1 == stateReg ? $signed(_GEN_393) : $signed({{16{_GEN_68[10]}},_GEN_68}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1433 = 3'h1 == stateReg ? $signed(_GEN_397) : $signed({{16{_GEN_70[10]}},_GEN_70}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1437 = 3'h1 == stateReg ? $signed(_GEN_401) : $signed({{16{_GEN_72[10]}},_GEN_72}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1441 = 3'h1 == stateReg ? $signed(_GEN_405) : $signed({{16{_GEN_74[10]}},_GEN_74}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1445 = 3'h1 == stateReg ? $signed(_GEN_409) : $signed({{16{_GEN_76[10]}},_GEN_76}); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire  _GEN_1544 = 3'h1 == stateReg ? 1'h0 : _GEN_1316; // @[\\src\\main\\scala\\GameLogic.scala 279:20 100:22]
  wire [26:0] _GEN_1548 = 3'h0 == stateReg ? $signed({{16{_GEN_18[10]}},_GEN_18}) : $signed(_GEN_1319); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1553 = 3'h0 == stateReg ? $signed({{16{_GEN_20[10]}},_GEN_20}) : $signed(_GEN_1324); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1558 = 3'h0 == stateReg ? $signed({{16{_GEN_22[10]}},_GEN_22}) : $signed(_GEN_1329); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1563 = 3'h0 == stateReg ? $signed({{16{_GEN_24[10]}},_GEN_24}) : $signed(_GEN_1334); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1568 = 3'h0 == stateReg ? $signed({{16{_GEN_26[10]}},_GEN_26}) : $signed(_GEN_1339); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1573 = 3'h0 == stateReg ? $signed({{16{_GEN_28[10]}},_GEN_28}) : $signed(_GEN_1344); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1578 = 3'h0 == stateReg ? $signed({{16{_GEN_30[10]}},_GEN_30}) : $signed(_GEN_1349); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1583 = 3'h0 == stateReg ? $signed({{16{_GEN_32[10]}},_GEN_32}) : $signed(_GEN_1354); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1588 = 3'h0 == stateReg ? $signed({{16{_GEN_34[10]}},_GEN_34}) : $signed(_GEN_1359); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1593 = 3'h0 == stateReg ? $signed({{16{_GEN_36[10]}},_GEN_36}) : $signed(_GEN_1364); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1598 = 3'h0 == stateReg ? $signed({{16{_GEN_38[10]}},_GEN_38}) : $signed(_GEN_1369); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1602 = 3'h0 == stateReg ? $signed({{16{_GEN_40[10]}},_GEN_40}) : $signed(_GEN_1373); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1606 = 3'h0 == stateReg ? $signed({{16{_GEN_42[10]}},_GEN_42}) : $signed(_GEN_1377); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1610 = 3'h0 == stateReg ? $signed({{16{_GEN_44[10]}},_GEN_44}) : $signed(_GEN_1381); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1614 = 3'h0 == stateReg ? $signed({{16{_GEN_46[10]}},_GEN_46}) : $signed(_GEN_1385); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1618 = 3'h0 == stateReg ? $signed({{16{_GEN_48[10]}},_GEN_48}) : $signed(_GEN_1389); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1622 = 3'h0 == stateReg ? $signed({{16{_GEN_50[10]}},_GEN_50}) : $signed(_GEN_1393); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1626 = 3'h0 == stateReg ? $signed({{16{_GEN_52[10]}},_GEN_52}) : $signed(_GEN_1397); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1630 = 3'h0 == stateReg ? $signed({{16{_GEN_54[10]}},_GEN_54}) : $signed(_GEN_1401); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1634 = 3'h0 == stateReg ? $signed({{16{_GEN_56[10]}},_GEN_56}) : $signed(_GEN_1405); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1638 = 3'h0 == stateReg ? $signed({{16{_GEN_58[10]}},_GEN_58}) : $signed(_GEN_1409); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1642 = 3'h0 == stateReg ? $signed({{16{_GEN_60[10]}},_GEN_60}) : $signed(_GEN_1413); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1646 = 3'h0 == stateReg ? $signed({{16{_GEN_62[10]}},_GEN_62}) : $signed(_GEN_1417); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1650 = 3'h0 == stateReg ? $signed({{16{_GEN_64[10]}},_GEN_64}) : $signed(_GEN_1421); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1654 = 3'h0 == stateReg ? $signed({{16{_GEN_66[10]}},_GEN_66}) : $signed(_GEN_1425); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1658 = 3'h0 == stateReg ? $signed({{16{_GEN_68[10]}},_GEN_68}) : $signed(_GEN_1429); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1662 = 3'h0 == stateReg ? $signed({{16{_GEN_70[10]}},_GEN_70}) : $signed(_GEN_1433); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1666 = 3'h0 == stateReg ? $signed({{16{_GEN_72[10]}},_GEN_72}) : $signed(_GEN_1437); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1670 = 3'h0 == stateReg ? $signed({{16{_GEN_74[10]}},_GEN_74}) : $signed(_GEN_1441); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1674 = 3'h0 == stateReg ? $signed({{16{_GEN_76[10]}},_GEN_76}) : $signed(_GEN_1445); // @[\\src\\main\\scala\\GameLogic.scala 279:20]
  wire [26:0] _GEN_1908 = reset ? $signed(27'sh0) : $signed(_GEN_1548); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1910 = reset ? $signed(27'sh0) : $signed(_GEN_1553); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1912 = reset ? $signed(27'sh0) : $signed(_GEN_1558); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1914 = reset ? $signed(27'sh0) : $signed(_GEN_1563); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1916 = reset ? $signed(27'sh0) : $signed(_GEN_1568); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1918 = reset ? $signed(27'sh0) : $signed(_GEN_1573); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1920 = reset ? $signed(27'sh0) : $signed(_GEN_1578); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1922 = reset ? $signed(27'sh0) : $signed(_GEN_1583); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1924 = reset ? $signed(27'sh0) : $signed(_GEN_1588); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1926 = reset ? $signed(27'sh0) : $signed(_GEN_1593); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1928 = reset ? $signed(27'sh0) : $signed(_GEN_1598); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1930 = reset ? $signed(27'sh0) : $signed(_GEN_1602); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1932 = reset ? $signed(27'sh0) : $signed(_GEN_1606); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1934 = reset ? $signed(27'sh0) : $signed(_GEN_1610); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1936 = reset ? $signed(27'sh0) : $signed(_GEN_1614); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1938 = reset ? $signed(27'sh0) : $signed(_GEN_1618); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1940 = reset ? $signed(27'sh0) : $signed(_GEN_1622); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1942 = reset ? $signed(27'sh0) : $signed(_GEN_1626); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1944 = reset ? $signed(27'sh0) : $signed(_GEN_1630); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1946 = reset ? $signed(27'sh0) : $signed(_GEN_1634); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1948 = reset ? $signed(27'sh0) : $signed(_GEN_1638); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1950 = reset ? $signed(27'sh0) : $signed(_GEN_1642); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1952 = reset ? $signed(27'sh0) : $signed(_GEN_1646); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1954 = reset ? $signed(27'sh0) : $signed(_GEN_1650); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1956 = reset ? $signed(27'sh0) : $signed(_GEN_1654); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1958 = reset ? $signed(27'sh0) : $signed(_GEN_1658); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1960 = reset ? $signed(27'sh0) : $signed(_GEN_1662); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1962 = reset ? $signed(27'sh0) : $signed(_GEN_1666); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1964 = reset ? $signed(27'sh0) : $signed(_GEN_1670); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_1966 = reset ? $signed(27'sh0) : $signed(_GEN_1674); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  Difficulty difficulty ( // @[\\src\\main\\scala\\GameLogic.scala 210:26]
    .clock(difficulty_clock),
    .reset(difficulty_reset),
    .io_level(difficulty_io_level),
    .io_speed(difficulty_io_speed),
    .io_resetSpeed(difficulty_io_resetSpeed)
  );
  LFSR lfsr ( // @[\\src\\main\\scala\\GameLogic.scala 248:20]
    .clock(lfsr_clock),
    .reset(lfsr_reset),
    .io_out_0(lfsr_io_out_0),
    .io_out_1(lfsr_io_out_1),
    .io_out_2(lfsr_io_out_2),
    .io_out_3(lfsr_io_out_3),
    .io_out_4(lfsr_io_out_4),
    .io_out_5(lfsr_io_out_5),
    .io_out_6(lfsr_io_out_6),
    .io_out_7(lfsr_io_out_7),
    .io_out_8(lfsr_io_out_8),
    .io_out_9(lfsr_io_out_9),
    .io_out_20(lfsr_io_out_20),
    .io_out_21(lfsr_io_out_21),
    .io_out_22(lfsr_io_out_22),
    .io_out_23(lfsr_io_out_23),
    .io_out_24(lfsr_io_out_24),
    .io_out_25(lfsr_io_out_25),
    .io_out_26(lfsr_io_out_26),
    .io_out_27(lfsr_io_out_27),
    .io_out_28(lfsr_io_out_28),
    .io_out_29(lfsr_io_out_29)
  );
  assign io_spriteXPosition_3 = spriteXRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_7 = spriteXRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_8 = spriteXRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_9 = spriteXRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_10 = spriteXRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_11 = spriteXRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_12 = spriteXRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_13 = spriteXRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_14 = spriteXRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_16 = spriteXRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_17 = spriteXRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_18 = spriteXRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_19 = spriteXRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_20 = spriteXRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_21 = spriteXRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_22 = spriteXRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_23 = spriteXRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_24 = spriteXRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_25 = spriteXRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_26 = spriteXRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_27 = spriteXRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_28 = spriteXRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_29 = spriteXRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_30 = spriteXRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_31 = spriteXRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_32 = spriteXRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_33 = spriteXRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_34 = spriteXRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_35 = spriteXRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_36 = spriteXRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_37 = spriteXRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_38 = spriteXRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_39 = spriteXRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_40 = spriteXRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_41 = spriteXRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_42 = spriteXRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_43 = spriteXRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_44 = spriteXRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_45 = spriteXRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_46 = spriteXRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_47 = spriteXRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_48 = spriteXRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_49 = spriteXRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_50 = spriteXRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_51 = spriteXRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_52 = spriteXRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_53 = spriteXRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_54 = spriteXRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_55 = spriteXRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_56 = spriteXRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_57 = spriteXRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_58 = spriteXRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_59 = spriteXRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_60 = spriteXRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_61 = spriteXRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_62 = spriteXRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteXPosition_63 = spriteXRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_3 = spriteYRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_7 = spriteYRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_8 = spriteYRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_9 = spriteYRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_10 = spriteYRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_11 = spriteYRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_12 = spriteYRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_13 = spriteYRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_14 = spriteYRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_16 = spriteYRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_17 = spriteYRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_18 = spriteYRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_19 = spriteYRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_20 = spriteYRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_21 = spriteYRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_22 = spriteYRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_23 = spriteYRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_24 = spriteYRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_25 = spriteYRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_26 = spriteYRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_27 = spriteYRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_28 = spriteYRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_29 = spriteYRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_30 = spriteYRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_31 = spriteYRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_32 = spriteYRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_33 = spriteYRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_34 = spriteYRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_35 = spriteYRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_36 = spriteYRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_37 = spriteYRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_38 = spriteYRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_39 = spriteYRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_40 = spriteYRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_41 = spriteYRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_42 = spriteYRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_43 = spriteYRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_44 = spriteYRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_45 = spriteYRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_46 = spriteYRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_47 = spriteYRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_48 = spriteYRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_49 = spriteYRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_50 = spriteYRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_51 = spriteYRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_52 = spriteYRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_53 = spriteYRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_54 = spriteYRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_55 = spriteYRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_56 = spriteYRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_57 = spriteYRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_58 = spriteYRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_59 = spriteYRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_60 = spriteYRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_61 = spriteYRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_62 = spriteYRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteYPosition_63 = spriteYRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 182:27]
  assign io_spriteVisible_3 = spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_4 = spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_5 = spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_6 = spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_7 = spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_8 = spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_9 = spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_10 = spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_11 = spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_12 = spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_13 = spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_14 = spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_15 = spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_16 = spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_17 = spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_18 = spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_19 = spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_20 = spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_21 = spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_22 = spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_23 = spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_24 = spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_25 = spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_26 = spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_27 = spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_28 = spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_29 = spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_30 = spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_31 = spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_32 = spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_33 = spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_34 = spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_35 = spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_36 = spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_37 = spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_38 = spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_39 = spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_40 = spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_41 = spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_42 = spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_43 = spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_44 = spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_45 = spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_46 = spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_47 = spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_48 = spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_49 = spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_50 = spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_51 = spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_52 = spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_53 = spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_54 = spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_55 = spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_56 = spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_57 = spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_58 = spriteVisibleRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_59 = spriteVisibleRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_60 = spriteVisibleRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_61 = spriteVisibleRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_62 = spriteVisibleRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteVisible_63 = spriteVisibleRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 178:25]
  assign io_spriteScaleUpHorizontal_16 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1322; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_17 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1327; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_18 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1332; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_19 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1337; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_20 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1342; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_21 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1347; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_22 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1352; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_23 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1357; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_24 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1362; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_25 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1367; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_26 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1322; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_27 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1327; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_28 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1332; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_29 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1337; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_30 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1342; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_31 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1347; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_32 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1352; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_33 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1357; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_34 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1362; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_35 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1367; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_36 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1322; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_37 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1327; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_38 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1332; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_39 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1337; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_40 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1342; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_41 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1347; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_42 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1352; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_43 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1357; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_44 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1362; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_45 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1367; // @[\\src\\main\\scala\\GameLogic.scala 279:20 188:33]
  assign io_spriteScaleUpHorizontal_58 = sprite58ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 194:34]
  assign io_spriteScaleUpHorizontal_59 = sprite59ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 196:34]
  assign io_spriteScaleUpHorizontal_60 = sprite60ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 198:34]
  assign io_spriteScaleUpVertical_16 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1322; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_17 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1327; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_18 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1332; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_19 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1337; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_20 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1342; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_21 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1347; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_22 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1352; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_23 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1357; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_24 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1362; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_25 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1367; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_26 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1322; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_27 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1327; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_28 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1332; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_29 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1337; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_30 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1342; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_31 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1347; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_32 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1352; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_33 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1357; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_34 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1362; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_35 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1367; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_36 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1322; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_37 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1327; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_38 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1332; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_39 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1337; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_40 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1342; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_41 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1347; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_42 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1352; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_43 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1357; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_44 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1362; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_45 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1367; // @[\\src\\main\\scala\\GameLogic.scala 279:20 189:31]
  assign io_spriteScaleUpVertical_58 = sprite58ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 195:32]
  assign io_spriteScaleUpVertical_59 = sprite59ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 197:32]
  assign io_spriteScaleUpVertical_60 = sprite60ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 199:32]
  assign io_viewBoxX = viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 206:15]
  assign io_viewBoxY = viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 207:15]
  assign io_frameUpdateDone = 3'h0 == stateReg ? 1'h0 : _GEN_1544; // @[\\src\\main\\scala\\GameLogic.scala 279:20 100:22]
  assign difficulty_clock = clock;
  assign difficulty_reset = reset;
  assign difficulty_io_level = lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 213:23]
  assign difficulty_io_resetSpeed = stateReg == 3'h2 & livesReg == 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 229:50]
  assign lfsr_clock = clock;
  assign lfsr_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 113:25]
      stateReg <= 3'h0; // @[\\src\\main\\scala\\GameLogic.scala 113:25]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 281:25]
        stateReg <= 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 282:18]
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (livesReg > 3'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 602:28]
        stateReg <= 3'h2; // @[\\src\\main\\scala\\GameLogic.scala 603:18]
      end else begin
        stateReg <= _GEN_1063;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      stateReg <= _GEN_1168;
    end else begin
      stateReg <= _GEN_1262;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_3 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_3 <= _GEN_0;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_3 <= _GEN_0;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_3 <= _GEN_0;
    end else begin
      spriteXRegs_3 <= _GEN_1264;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_7 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_7 <= 11'sh100; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_8 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_8 <= 11'sh100; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_9 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_9 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_10 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_10 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_11 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_11 <= 11'sh160; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_12 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_12 <= 11'sh160; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_13 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_13 <= _GEN_14;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteXRegs_13 <= _GEN_281;
      end else begin
        spriteXRegs_13 <= _GEN_14;
      end
    end else begin
      spriteXRegs_13 <= _GEN_14;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_14 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_14 <= _GEN_16;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_14 <= _GEN_16;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_14 <= _GEN_16;
    end else begin
      spriteXRegs_14 <= _GEN_1247;
    end
    spriteXRegs_16 <= _GEN_1908[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_17 <= _GEN_1910[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_18 <= _GEN_1912[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_19 <= _GEN_1914[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_20 <= _GEN_1916[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_21 <= _GEN_1918[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_22 <= _GEN_1920[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_23 <= _GEN_1922[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_24 <= _GEN_1924[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_25 <= _GEN_1926[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_26 <= _GEN_1928[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_27 <= _GEN_1930[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_28 <= _GEN_1932[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_29 <= _GEN_1934[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_30 <= _GEN_1936[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_31 <= _GEN_1938[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_32 <= _GEN_1940[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_33 <= _GEN_1942[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_34 <= _GEN_1944[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_35 <= _GEN_1946[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_36 <= _GEN_1948[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_37 <= _GEN_1950[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_38 <= _GEN_1952[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_39 <= _GEN_1954[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_40 <= _GEN_1956[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_41 <= _GEN_1958[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_42 <= _GEN_1960[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_43 <= _GEN_1962[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_44 <= _GEN_1964[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_45 <= _GEN_1966[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_46 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_46 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_47 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_47 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_48 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_48 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_49 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_49 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_50 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_50 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_51 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_51 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_52 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_52 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_53 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_53 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_54 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_54 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_55 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_55 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_56 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_56 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_57 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_57 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_58 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_58 <= _GEN_102;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 512:29]
        spriteXRegs_58 <= spriteXRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 513:25]
      end else begin
        spriteXRegs_58 <= _GEN_1125;
      end
    end else begin
      spriteXRegs_58 <= _GEN_102;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_59 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_59 <= _GEN_104;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 512:29]
        spriteXRegs_59 <= spriteXRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 515:25]
      end else begin
        spriteXRegs_59 <= _GEN_1126;
      end
    end else begin
      spriteXRegs_59 <= _GEN_104;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_60 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteXRegs_60 <= _GEN_106;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 512:29]
        spriteXRegs_60 <= spriteXRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 517:25]
      end else begin
        spriteXRegs_60 <= _GEN_1127;
      end
    end else begin
      spriteXRegs_60 <= _GEN_106;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_61 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_61 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_62 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_62 <= 11'sh3c; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_63 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteXRegs_63 <= 11'sh64; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_3 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_3 <= _GEN_1;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_3 <= _GEN_1;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_3 <= _GEN_1;
    end else begin
      spriteYRegs_3 <= _GEN_1263;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_7 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_7 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_8 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_8 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_9 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_9 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_10 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_10 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_11 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_11 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_12 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_12 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_13 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_13 <= _GEN_15;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_13 <= _GEN_279;
      end else begin
        spriteYRegs_13 <= _GEN_15;
      end
    end else begin
      spriteYRegs_13 <= _GEN_15;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_14 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_14 <= _GEN_17;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_14 <= _GEN_17;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_14 <= _GEN_17;
    end else begin
      spriteYRegs_14 <= _GEN_1248;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_16 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_16 <= _GEN_19;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_16 <= _GEN_129;
      end else begin
        spriteYRegs_16 <= _GEN_19;
      end
    end else begin
      spriteYRegs_16 <= _GEN_19;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_17 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_17 <= _GEN_21;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_17 <= _GEN_134;
      end else begin
        spriteYRegs_17 <= _GEN_21;
      end
    end else begin
      spriteYRegs_17 <= _GEN_21;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_18 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_18 <= _GEN_23;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_18 <= _GEN_139;
      end else begin
        spriteYRegs_18 <= _GEN_23;
      end
    end else begin
      spriteYRegs_18 <= _GEN_23;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_19 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_19 <= _GEN_25;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_19 <= _GEN_144;
      end else begin
        spriteYRegs_19 <= _GEN_25;
      end
    end else begin
      spriteYRegs_19 <= _GEN_25;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_20 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_20 <= _GEN_27;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_20 <= _GEN_149;
      end else begin
        spriteYRegs_20 <= _GEN_27;
      end
    end else begin
      spriteYRegs_20 <= _GEN_27;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_21 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_21 <= _GEN_29;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_21 <= _GEN_154;
      end else begin
        spriteYRegs_21 <= _GEN_29;
      end
    end else begin
      spriteYRegs_21 <= _GEN_29;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_22 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_22 <= _GEN_31;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_22 <= _GEN_159;
      end else begin
        spriteYRegs_22 <= _GEN_31;
      end
    end else begin
      spriteYRegs_22 <= _GEN_31;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_23 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_23 <= _GEN_33;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_23 <= _GEN_164;
      end else begin
        spriteYRegs_23 <= _GEN_33;
      end
    end else begin
      spriteYRegs_23 <= _GEN_33;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_24 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_24 <= _GEN_35;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_24 <= _GEN_169;
      end else begin
        spriteYRegs_24 <= _GEN_35;
      end
    end else begin
      spriteYRegs_24 <= _GEN_35;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_25 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_25 <= _GEN_37;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_25 <= _GEN_174;
      end else begin
        spriteYRegs_25 <= _GEN_37;
      end
    end else begin
      spriteYRegs_25 <= _GEN_37;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_26 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_26 <= _GEN_39;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_26 <= _GEN_179;
      end else begin
        spriteYRegs_26 <= _GEN_39;
      end
    end else begin
      spriteYRegs_26 <= _GEN_39;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_27 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_27 <= _GEN_41;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_27 <= _GEN_184;
      end else begin
        spriteYRegs_27 <= _GEN_41;
      end
    end else begin
      spriteYRegs_27 <= _GEN_41;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_28 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_28 <= _GEN_43;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_28 <= _GEN_189;
      end else begin
        spriteYRegs_28 <= _GEN_43;
      end
    end else begin
      spriteYRegs_28 <= _GEN_43;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_29 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_29 <= _GEN_45;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_29 <= _GEN_194;
      end else begin
        spriteYRegs_29 <= _GEN_45;
      end
    end else begin
      spriteYRegs_29 <= _GEN_45;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_30 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_30 <= _GEN_47;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_30 <= _GEN_199;
      end else begin
        spriteYRegs_30 <= _GEN_47;
      end
    end else begin
      spriteYRegs_30 <= _GEN_47;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_31 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_31 <= _GEN_49;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_31 <= _GEN_204;
      end else begin
        spriteYRegs_31 <= _GEN_49;
      end
    end else begin
      spriteYRegs_31 <= _GEN_49;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_32 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_32 <= _GEN_51;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_32 <= _GEN_209;
      end else begin
        spriteYRegs_32 <= _GEN_51;
      end
    end else begin
      spriteYRegs_32 <= _GEN_51;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_33 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_33 <= _GEN_53;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_33 <= _GEN_214;
      end else begin
        spriteYRegs_33 <= _GEN_53;
      end
    end else begin
      spriteYRegs_33 <= _GEN_53;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_34 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_34 <= _GEN_55;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_34 <= _GEN_219;
      end else begin
        spriteYRegs_34 <= _GEN_55;
      end
    end else begin
      spriteYRegs_34 <= _GEN_55;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_35 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_35 <= _GEN_57;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_35 <= _GEN_224;
      end else begin
        spriteYRegs_35 <= _GEN_57;
      end
    end else begin
      spriteYRegs_35 <= _GEN_57;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_36 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_36 <= _GEN_59;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_36 <= _GEN_229;
      end else begin
        spriteYRegs_36 <= _GEN_59;
      end
    end else begin
      spriteYRegs_36 <= _GEN_59;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_37 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_37 <= _GEN_61;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_37 <= _GEN_234;
      end else begin
        spriteYRegs_37 <= _GEN_61;
      end
    end else begin
      spriteYRegs_37 <= _GEN_61;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_38 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_38 <= _GEN_63;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_38 <= _GEN_239;
      end else begin
        spriteYRegs_38 <= _GEN_63;
      end
    end else begin
      spriteYRegs_38 <= _GEN_63;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_39 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_39 <= _GEN_65;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_39 <= _GEN_244;
      end else begin
        spriteYRegs_39 <= _GEN_65;
      end
    end else begin
      spriteYRegs_39 <= _GEN_65;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_40 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_40 <= _GEN_67;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_40 <= _GEN_249;
      end else begin
        spriteYRegs_40 <= _GEN_67;
      end
    end else begin
      spriteYRegs_40 <= _GEN_67;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_41 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_41 <= _GEN_69;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_41 <= _GEN_254;
      end else begin
        spriteYRegs_41 <= _GEN_69;
      end
    end else begin
      spriteYRegs_41 <= _GEN_69;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_42 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_42 <= _GEN_71;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_42 <= _GEN_259;
      end else begin
        spriteYRegs_42 <= _GEN_71;
      end
    end else begin
      spriteYRegs_42 <= _GEN_71;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_43 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_43 <= _GEN_73;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_43 <= _GEN_264;
      end else begin
        spriteYRegs_43 <= _GEN_73;
      end
    end else begin
      spriteYRegs_43 <= _GEN_73;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_44 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_44 <= _GEN_75;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_44 <= _GEN_269;
      end else begin
        spriteYRegs_44 <= _GEN_75;
      end
    end else begin
      spriteYRegs_44 <= _GEN_75;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_45 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_45 <= _GEN_77;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
        spriteYRegs_45 <= _GEN_274;
      end else begin
        spriteYRegs_45 <= _GEN_77;
      end
    end else begin
      spriteYRegs_45 <= _GEN_77;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_46 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_46 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_47 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_47 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_48 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_48 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_49 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_49 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_50 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_50 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_51 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_51 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_52 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_52 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_53 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_53 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_54 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_54 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_55 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_55 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_56 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_56 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_57 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_57 <= 10'sh122; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_58 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_58 <= _GEN_103;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 512:29]
        spriteYRegs_58 <= spriteYRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 514:25]
      end else begin
        spriteYRegs_58 <= _GEN_1128;
      end
    end else begin
      spriteYRegs_58 <= _GEN_103;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_59 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_59 <= _GEN_105;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 512:29]
        spriteYRegs_59 <= spriteYRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 516:25]
      end else begin
        spriteYRegs_59 <= _GEN_1129;
      end
    end else begin
      spriteYRegs_59 <= _GEN_105;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_60 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteYRegs_60 <= _GEN_107;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 512:29]
        spriteYRegs_60 <= spriteYRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 518:25]
      end else begin
        spriteYRegs_60 <= _GEN_1130;
      end
    end else begin
      spriteYRegs_60 <= _GEN_107;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_61 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_61 <= 10'sh14; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_62 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_62 <= 10'sh14; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_63 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 132:29]
      spriteYRegs_63 <= 10'sh14; // @[\\src\\main\\scala\\GameLogic.scala 163:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_3 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_3 <= _GEN_485;
        end else begin
          spriteVisibleRegs_3 <= _GEN_879;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_3 <= _GEN_1169;
      end else begin
        spriteVisibleRegs_3 <= _GEN_1249;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_4 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_4 <= _GEN_486;
        end else begin
          spriteVisibleRegs_4 <= _GEN_880;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_5 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_5 <= _GEN_487;
        end else begin
          spriteVisibleRegs_5 <= _GEN_881;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_6 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_6 <= _GEN_488;
        end else begin
          spriteVisibleRegs_6 <= _GEN_882;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_7 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_7 <= _GEN_489;
        end else begin
          spriteVisibleRegs_7 <= _GEN_883;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_7 <= _GEN_1170;
      end else begin
        spriteVisibleRegs_7 <= _GEN_1250;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_8 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_8 <= _GEN_490;
        end else begin
          spriteVisibleRegs_8 <= _GEN_884;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_8 <= _GEN_1171;
      end else begin
        spriteVisibleRegs_8 <= _GEN_1251;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_9 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_9 <= _GEN_491;
        end else begin
          spriteVisibleRegs_9 <= _GEN_885;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_9 <= _GEN_1172;
      end else begin
        spriteVisibleRegs_9 <= _GEN_1252;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_10 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_10 <= _GEN_492;
        end else begin
          spriteVisibleRegs_10 <= _GEN_886;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_10 <= _GEN_1173;
      end else begin
        spriteVisibleRegs_10 <= _GEN_1253;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_11 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_11 <= _GEN_493;
        end else begin
          spriteVisibleRegs_11 <= _GEN_887;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_11 <= _GEN_1174;
      end else begin
        spriteVisibleRegs_11 <= _GEN_1254;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_12 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_12 <= _GEN_494;
        end else begin
          spriteVisibleRegs_12 <= _GEN_888;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_12 <= _GEN_1175;
      end else begin
        spriteVisibleRegs_12 <= _GEN_1255;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_13 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T_731) begin // @[\\src\\main\\scala\\GameLogic.scala 458:9]
          spriteVisibleRegs_13 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 459:31]
        end else begin
          spriteVisibleRegs_13 <= _GEN_955;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_14 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 473:24]
          spriteVisibleRegs_14 <= _GEN_1054;
        end else begin
          spriteVisibleRegs_14 <= _GEN_956;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_14 <= _GEN_1256;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_15 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_15 <= _GEN_497;
        end else begin
          spriteVisibleRegs_15 <= _GEN_891;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_16 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_16 <= _GEN_498;
        end else begin
          spriteVisibleRegs_16 <= _GEN_892;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_17 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_17 <= _GEN_499;
        end else begin
          spriteVisibleRegs_17 <= _GEN_893;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_18 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_18 <= _GEN_500;
        end else begin
          spriteVisibleRegs_18 <= _GEN_894;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_19 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_19 <= _GEN_501;
        end else begin
          spriteVisibleRegs_19 <= _GEN_895;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_20 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_20 <= _GEN_502;
        end else begin
          spriteVisibleRegs_20 <= _GEN_896;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_21 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_21 <= _GEN_503;
        end else begin
          spriteVisibleRegs_21 <= _GEN_897;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_22 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_22 <= _GEN_504;
        end else begin
          spriteVisibleRegs_22 <= _GEN_898;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_23 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_23 <= _GEN_505;
        end else begin
          spriteVisibleRegs_23 <= _GEN_899;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_24 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_24 <= _GEN_506;
        end else begin
          spriteVisibleRegs_24 <= _GEN_900;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_25 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_25 <= _GEN_507;
        end else begin
          spriteVisibleRegs_25 <= _GEN_901;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_26 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_26 <= _GEN_508;
        end else begin
          spriteVisibleRegs_26 <= _GEN_902;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_27 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_27 <= _GEN_509;
        end else begin
          spriteVisibleRegs_27 <= _GEN_903;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_28 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_28 <= _GEN_510;
        end else begin
          spriteVisibleRegs_28 <= _GEN_904;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_29 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_29 <= _GEN_511;
        end else begin
          spriteVisibleRegs_29 <= _GEN_905;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_30 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_30 <= _GEN_512;
        end else begin
          spriteVisibleRegs_30 <= _GEN_906;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_31 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_31 <= _GEN_513;
        end else begin
          spriteVisibleRegs_31 <= _GEN_907;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_32 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_32 <= _GEN_514;
        end else begin
          spriteVisibleRegs_32 <= _GEN_908;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_33 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_33 <= _GEN_515;
        end else begin
          spriteVisibleRegs_33 <= _GEN_909;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_34 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_34 <= _GEN_516;
        end else begin
          spriteVisibleRegs_34 <= _GEN_910;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_35 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_35 <= _GEN_517;
        end else begin
          spriteVisibleRegs_35 <= _GEN_911;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_36 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_36 <= _GEN_518;
        end else begin
          spriteVisibleRegs_36 <= _GEN_912;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_37 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_37 <= _GEN_519;
        end else begin
          spriteVisibleRegs_37 <= _GEN_913;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_38 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_38 <= _GEN_520;
        end else begin
          spriteVisibleRegs_38 <= _GEN_914;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_39 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_39 <= _GEN_521;
        end else begin
          spriteVisibleRegs_39 <= _GEN_915;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_40 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_40 <= _GEN_522;
        end else begin
          spriteVisibleRegs_40 <= _GEN_916;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_41 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_41 <= _GEN_523;
        end else begin
          spriteVisibleRegs_41 <= _GEN_917;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_42 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_42 <= _GEN_524;
        end else begin
          spriteVisibleRegs_42 <= _GEN_918;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_43 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_43 <= _GEN_525;
        end else begin
          spriteVisibleRegs_43 <= _GEN_919;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_44 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_44 <= _GEN_526;
        end else begin
          spriteVisibleRegs_44 <= _GEN_920;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_45 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_45 <= _GEN_527;
        end else begin
          spriteVisibleRegs_45 <= _GEN_921;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_46 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_46 <= _GEN_528;
        end else begin
          spriteVisibleRegs_46 <= _GEN_922;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_46 <= _GEN_1265;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_47 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_47 <= _GEN_529;
        end else begin
          spriteVisibleRegs_47 <= _GEN_923;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_47 <= _GEN_1266;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_48 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_48 <= _GEN_530;
        end else begin
          spriteVisibleRegs_48 <= _GEN_924;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_48 <= _GEN_1267;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_49 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_49 <= _GEN_531;
        end else begin
          spriteVisibleRegs_49 <= _GEN_925;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_49 <= _GEN_1268;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_50 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_50 <= _GEN_532;
        end else begin
          spriteVisibleRegs_50 <= _GEN_926;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_50 <= _GEN_1269;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_51 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_51 <= _GEN_533;
        end else begin
          spriteVisibleRegs_51 <= _GEN_927;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_51 <= _GEN_1270;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_52 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_52 <= _GEN_534;
        end else begin
          spriteVisibleRegs_52 <= _GEN_928;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_52 <= _GEN_1271;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_53 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_53 <= _GEN_535;
        end else begin
          spriteVisibleRegs_53 <= _GEN_929;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_53 <= _GEN_1272;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_54 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_54 <= _GEN_536;
        end else begin
          spriteVisibleRegs_54 <= _GEN_930;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_54 <= _GEN_1273;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_55 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_55 <= _GEN_537;
        end else begin
          spriteVisibleRegs_55 <= _GEN_931;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_55 <= _GEN_1274;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_56 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_56 <= _GEN_538;
        end else begin
          spriteVisibleRegs_56 <= _GEN_932;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_56 <= _GEN_1275;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_57 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spriteVisibleRegs_57 <= _GEN_539;
        end else begin
          spriteVisibleRegs_57 <= _GEN_933;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_57 <= _GEN_1276;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_58 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_58 <= _T_82;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_59 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_59 <= _T_82;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_60 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spriteVisibleRegs_60 <= _T_82;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_61 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteVisibleRegs_61 <= _GEN_123;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
        spriteVisibleRegs_61 <= _GEN_543;
      end else begin
        spriteVisibleRegs_61 <= _GEN_937;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteVisibleRegs_61 <= _GEN_123;
    end else begin
      spriteVisibleRegs_61 <= _GEN_1257;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_62 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteVisibleRegs_62 <= _GEN_124;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
        spriteVisibleRegs_62 <= _GEN_544;
      end else begin
        spriteVisibleRegs_62 <= _GEN_938;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteVisibleRegs_62 <= _GEN_124;
    end else begin
      spriteVisibleRegs_62 <= _GEN_1258;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_63 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteVisibleRegs_63 <= _GEN_125;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
        spriteVisibleRegs_63 <= _GEN_545;
      end else begin
        spriteVisibleRegs_63 <= _GEN_939;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      spriteVisibleRegs_63 <= _GEN_125;
    end else begin
      spriteVisibleRegs_63 <= _GEN_1259;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_0 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_0 <= _GEN_230;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_1 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_1 <= _GEN_235;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_2 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_2 <= _GEN_240;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_3 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_3 <= _GEN_245;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_4 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_4 <= _GEN_250;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_5 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_5 <= _GEN_255;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_6 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_6 <= _GEN_260;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_7 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_7 <= _GEN_265;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_8 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_8 <= _GEN_270;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_9 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          spriteScaleTypeRegs_9 <= _GEN_275;
        end
      end
    end
    initializePositions <= reset | _GEN_114; // @[\\src\\main\\scala\\GameLogic.scala 131:{36,36}]
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 169:42]
      sprite58ScaleUpHorizontal <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 169:42]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        sprite58ScaleUpHorizontal <= _GEN_1138;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 170:40]
      sprite58ScaleUpVertical <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 170:40]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        sprite58ScaleUpVertical <= _GEN_1141;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 171:42]
      sprite59ScaleUpHorizontal <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 171:42]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        sprite59ScaleUpHorizontal <= _GEN_1139;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 172:40]
      sprite59ScaleUpVertical <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 172:40]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        sprite59ScaleUpVertical <= _GEN_1142;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 173:42]
      sprite60ScaleUpHorizontal <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 173:42]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        sprite60ScaleUpHorizontal <= _GEN_1140;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 174:40]
      sprite60ScaleUpVertical <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 174:40]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        sprite60ScaleUpVertical <= _GEN_1143;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 202:28]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 202:28]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
          viewBoxXReg <= _GEN_1260;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 203:28]
      viewBoxYReg <= 9'h0; // @[\\src\\main\\scala\\GameLogic.scala 203:28]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
          viewBoxYReg <= _GEN_1261;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 212:23]
      lvlReg <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 212:23]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
          lvlReg <= _GEN_1176;
        end else begin
          lvlReg <= _GEN_1277;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 223:25]
      livesReg <= 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 223:25]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 473:24]
          livesReg <= _GEN_1055;
        end else begin
          livesReg <= _GEN_1043;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        livesReg <= _GEN_1278;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 226:29]
      extraLifeCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 226:29]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 294:29]
          extraLifeCnt <= _GEN_280;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 232:34]
      spawnDelayCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 232:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          spawnDelayCounter <= _GEN_547;
        end else begin
          spawnDelayCounter <= _GEN_941;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        spawnDelayCounter <= _GEN_1246;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 233:34]
      nextSpriteToSpawn <= 6'h0; // @[\\src\\main\\scala\\GameLogic.scala 233:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 385:28]
          nextSpriteToSpawn <= _GEN_546;
        end else begin
          nextSpriteToSpawn <= _GEN_940;
        end
      end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        nextSpriteToSpawn <= _GEN_1245;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 236:24]
      starCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 236:24]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 512:29]
          starCnt <= _starCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 525:17]
        end else begin
          starCnt <= _GEN_1131;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 239:34]
      collisionDetected <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 239:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 473:24]
          collisionDetected <= _GEN_1057;
        end else begin
          collisionDetected <= _GEN_1040;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 240:29]
      blinkCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 240:29]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 473:24]
          blinkCounter <= _GEN_1049;
        end else begin
          blinkCounter <= _GEN_1045;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 241:27]
      blinkTimes <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 241:27]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 473:24]
          blinkTimes <= _GEN_1050;
        end else begin
          blinkTimes <= _GEN_1046;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 242:27]
      isBlinking <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 242:27]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 279:20]
        if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 473:24]
          isBlinking <= _GEN_1053;
        end else begin
          isBlinking <= _GEN_1044;
        end
      end
    end
    spriteXRegs_58_REG <= $signed(spriteXRegs_59) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 513:52]
    spriteYRegs_58_REG <= $signed(spriteYRegs_59) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 514:52]
    spriteXRegs_59_REG <= $signed(spriteXRegs_60) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 515:52]
    spriteYRegs_59_REG <= $signed(spriteYRegs_60) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 516:52]
    spriteXRegs_60_REG <= $signed(spriteXRegs_58) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 517:52]
    spriteYRegs_60_REG <= $signed(spriteYRegs_58) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 518:52]
    spriteXRegs_58_REG_1 <= $signed(spriteXRegs_59) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 541:52]
    spriteYRegs_58_REG_1 <= $signed(spriteYRegs_59) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 542:52]
    spriteXRegs_59_REG_1 <= $signed(spriteXRegs_60) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 543:52]
    spriteYRegs_59_REG_1 <= $signed(spriteYRegs_60) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 544:52]
    spriteXRegs_60_REG_1 <= $signed(spriteXRegs_58) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 545:52]
    spriteYRegs_60_REG_1 <= $signed(spriteYRegs_58) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 546:52]
    spriteXRegs_58_REG_2 <= $signed(spriteXRegs_59) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 569:52]
    spriteYRegs_58_REG_2 <= $signed(spriteYRegs_59) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 570:52]
    spriteXRegs_59_REG_2 <= $signed(spriteXRegs_60) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 571:52]
    spriteYRegs_59_REG_2 <= $signed(spriteYRegs_60) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 572:52]
    spriteXRegs_60_REG_2 <= $signed(spriteXRegs_58) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 573:52]
    spriteYRegs_60_REG_2 <= $signed(spriteYRegs_58) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 574:52]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  spriteXRegs_3 = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  spriteXRegs_7 = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  spriteXRegs_8 = _RAND_3[10:0];
  _RAND_4 = {1{`RANDOM}};
  spriteXRegs_9 = _RAND_4[10:0];
  _RAND_5 = {1{`RANDOM}};
  spriteXRegs_10 = _RAND_5[10:0];
  _RAND_6 = {1{`RANDOM}};
  spriteXRegs_11 = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  spriteXRegs_12 = _RAND_7[10:0];
  _RAND_8 = {1{`RANDOM}};
  spriteXRegs_13 = _RAND_8[10:0];
  _RAND_9 = {1{`RANDOM}};
  spriteXRegs_14 = _RAND_9[10:0];
  _RAND_10 = {1{`RANDOM}};
  spriteXRegs_16 = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  spriteXRegs_17 = _RAND_11[10:0];
  _RAND_12 = {1{`RANDOM}};
  spriteXRegs_18 = _RAND_12[10:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXRegs_19 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXRegs_20 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXRegs_21 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXRegs_22 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXRegs_23 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXRegs_24 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXRegs_25 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteXRegs_26 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  spriteXRegs_27 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  spriteXRegs_28 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  spriteXRegs_29 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  spriteXRegs_30 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  spriteXRegs_31 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  spriteXRegs_32 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  spriteXRegs_33 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  spriteXRegs_34 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  spriteXRegs_35 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  spriteXRegs_36 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  spriteXRegs_37 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  spriteXRegs_38 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  spriteXRegs_39 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  spriteXRegs_40 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  spriteXRegs_41 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  spriteXRegs_42 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  spriteXRegs_43 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  spriteXRegs_44 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  spriteXRegs_45 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  spriteXRegs_46 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  spriteXRegs_47 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  spriteXRegs_48 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  spriteXRegs_49 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  spriteXRegs_50 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  spriteXRegs_51 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  spriteXRegs_52 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  spriteXRegs_53 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  spriteXRegs_54 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  spriteXRegs_55 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  spriteXRegs_56 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  spriteXRegs_57 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  spriteXRegs_58 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  spriteXRegs_59 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  spriteXRegs_60 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  spriteXRegs_61 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  spriteXRegs_62 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  spriteXRegs_63 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  spriteYRegs_3 = _RAND_58[9:0];
  _RAND_59 = {1{`RANDOM}};
  spriteYRegs_7 = _RAND_59[9:0];
  _RAND_60 = {1{`RANDOM}};
  spriteYRegs_8 = _RAND_60[9:0];
  _RAND_61 = {1{`RANDOM}};
  spriteYRegs_9 = _RAND_61[9:0];
  _RAND_62 = {1{`RANDOM}};
  spriteYRegs_10 = _RAND_62[9:0];
  _RAND_63 = {1{`RANDOM}};
  spriteYRegs_11 = _RAND_63[9:0];
  _RAND_64 = {1{`RANDOM}};
  spriteYRegs_12 = _RAND_64[9:0];
  _RAND_65 = {1{`RANDOM}};
  spriteYRegs_13 = _RAND_65[9:0];
  _RAND_66 = {1{`RANDOM}};
  spriteYRegs_14 = _RAND_66[9:0];
  _RAND_67 = {1{`RANDOM}};
  spriteYRegs_16 = _RAND_67[9:0];
  _RAND_68 = {1{`RANDOM}};
  spriteYRegs_17 = _RAND_68[9:0];
  _RAND_69 = {1{`RANDOM}};
  spriteYRegs_18 = _RAND_69[9:0];
  _RAND_70 = {1{`RANDOM}};
  spriteYRegs_19 = _RAND_70[9:0];
  _RAND_71 = {1{`RANDOM}};
  spriteYRegs_20 = _RAND_71[9:0];
  _RAND_72 = {1{`RANDOM}};
  spriteYRegs_21 = _RAND_72[9:0];
  _RAND_73 = {1{`RANDOM}};
  spriteYRegs_22 = _RAND_73[9:0];
  _RAND_74 = {1{`RANDOM}};
  spriteYRegs_23 = _RAND_74[9:0];
  _RAND_75 = {1{`RANDOM}};
  spriteYRegs_24 = _RAND_75[9:0];
  _RAND_76 = {1{`RANDOM}};
  spriteYRegs_25 = _RAND_76[9:0];
  _RAND_77 = {1{`RANDOM}};
  spriteYRegs_26 = _RAND_77[9:0];
  _RAND_78 = {1{`RANDOM}};
  spriteYRegs_27 = _RAND_78[9:0];
  _RAND_79 = {1{`RANDOM}};
  spriteYRegs_28 = _RAND_79[9:0];
  _RAND_80 = {1{`RANDOM}};
  spriteYRegs_29 = _RAND_80[9:0];
  _RAND_81 = {1{`RANDOM}};
  spriteYRegs_30 = _RAND_81[9:0];
  _RAND_82 = {1{`RANDOM}};
  spriteYRegs_31 = _RAND_82[9:0];
  _RAND_83 = {1{`RANDOM}};
  spriteYRegs_32 = _RAND_83[9:0];
  _RAND_84 = {1{`RANDOM}};
  spriteYRegs_33 = _RAND_84[9:0];
  _RAND_85 = {1{`RANDOM}};
  spriteYRegs_34 = _RAND_85[9:0];
  _RAND_86 = {1{`RANDOM}};
  spriteYRegs_35 = _RAND_86[9:0];
  _RAND_87 = {1{`RANDOM}};
  spriteYRegs_36 = _RAND_87[9:0];
  _RAND_88 = {1{`RANDOM}};
  spriteYRegs_37 = _RAND_88[9:0];
  _RAND_89 = {1{`RANDOM}};
  spriteYRegs_38 = _RAND_89[9:0];
  _RAND_90 = {1{`RANDOM}};
  spriteYRegs_39 = _RAND_90[9:0];
  _RAND_91 = {1{`RANDOM}};
  spriteYRegs_40 = _RAND_91[9:0];
  _RAND_92 = {1{`RANDOM}};
  spriteYRegs_41 = _RAND_92[9:0];
  _RAND_93 = {1{`RANDOM}};
  spriteYRegs_42 = _RAND_93[9:0];
  _RAND_94 = {1{`RANDOM}};
  spriteYRegs_43 = _RAND_94[9:0];
  _RAND_95 = {1{`RANDOM}};
  spriteYRegs_44 = _RAND_95[9:0];
  _RAND_96 = {1{`RANDOM}};
  spriteYRegs_45 = _RAND_96[9:0];
  _RAND_97 = {1{`RANDOM}};
  spriteYRegs_46 = _RAND_97[9:0];
  _RAND_98 = {1{`RANDOM}};
  spriteYRegs_47 = _RAND_98[9:0];
  _RAND_99 = {1{`RANDOM}};
  spriteYRegs_48 = _RAND_99[9:0];
  _RAND_100 = {1{`RANDOM}};
  spriteYRegs_49 = _RAND_100[9:0];
  _RAND_101 = {1{`RANDOM}};
  spriteYRegs_50 = _RAND_101[9:0];
  _RAND_102 = {1{`RANDOM}};
  spriteYRegs_51 = _RAND_102[9:0];
  _RAND_103 = {1{`RANDOM}};
  spriteYRegs_52 = _RAND_103[9:0];
  _RAND_104 = {1{`RANDOM}};
  spriteYRegs_53 = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  spriteYRegs_54 = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  spriteYRegs_55 = _RAND_106[9:0];
  _RAND_107 = {1{`RANDOM}};
  spriteYRegs_56 = _RAND_107[9:0];
  _RAND_108 = {1{`RANDOM}};
  spriteYRegs_57 = _RAND_108[9:0];
  _RAND_109 = {1{`RANDOM}};
  spriteYRegs_58 = _RAND_109[9:0];
  _RAND_110 = {1{`RANDOM}};
  spriteYRegs_59 = _RAND_110[9:0];
  _RAND_111 = {1{`RANDOM}};
  spriteYRegs_60 = _RAND_111[9:0];
  _RAND_112 = {1{`RANDOM}};
  spriteYRegs_61 = _RAND_112[9:0];
  _RAND_113 = {1{`RANDOM}};
  spriteYRegs_62 = _RAND_113[9:0];
  _RAND_114 = {1{`RANDOM}};
  spriteYRegs_63 = _RAND_114[9:0];
  _RAND_115 = {1{`RANDOM}};
  spriteVisibleRegs_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  spriteVisibleRegs_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  spriteVisibleRegs_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  spriteVisibleRegs_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  spriteVisibleRegs_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  spriteVisibleRegs_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  spriteVisibleRegs_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  spriteVisibleRegs_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  spriteVisibleRegs_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  spriteVisibleRegs_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  spriteVisibleRegs_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  spriteVisibleRegs_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  spriteVisibleRegs_15 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  spriteVisibleRegs_16 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  spriteVisibleRegs_17 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  spriteVisibleRegs_18 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  spriteVisibleRegs_19 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  spriteVisibleRegs_20 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  spriteVisibleRegs_21 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  spriteVisibleRegs_22 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  spriteVisibleRegs_23 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  spriteVisibleRegs_24 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  spriteVisibleRegs_25 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  spriteVisibleRegs_26 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  spriteVisibleRegs_27 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  spriteVisibleRegs_28 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  spriteVisibleRegs_29 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  spriteVisibleRegs_30 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  spriteVisibleRegs_31 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  spriteVisibleRegs_32 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  spriteVisibleRegs_33 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  spriteVisibleRegs_34 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  spriteVisibleRegs_35 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  spriteVisibleRegs_36 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  spriteVisibleRegs_37 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  spriteVisibleRegs_38 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  spriteVisibleRegs_39 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  spriteVisibleRegs_40 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  spriteVisibleRegs_41 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  spriteVisibleRegs_42 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  spriteVisibleRegs_43 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  spriteVisibleRegs_44 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  spriteVisibleRegs_45 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  spriteVisibleRegs_46 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  spriteVisibleRegs_47 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  spriteVisibleRegs_48 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  spriteVisibleRegs_49 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  spriteVisibleRegs_50 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  spriteVisibleRegs_51 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  spriteVisibleRegs_52 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  spriteVisibleRegs_53 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  spriteVisibleRegs_54 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  spriteVisibleRegs_55 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  spriteVisibleRegs_56 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  spriteVisibleRegs_57 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  spriteVisibleRegs_58 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  spriteVisibleRegs_59 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  spriteVisibleRegs_60 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  spriteVisibleRegs_61 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  spriteVisibleRegs_62 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  spriteVisibleRegs_63 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  spriteScaleTypeRegs_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  spriteScaleTypeRegs_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  spriteScaleTypeRegs_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  spriteScaleTypeRegs_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  spriteScaleTypeRegs_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  spriteScaleTypeRegs_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  spriteScaleTypeRegs_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  spriteScaleTypeRegs_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  spriteScaleTypeRegs_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  spriteScaleTypeRegs_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  initializePositions = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  sprite58ScaleUpHorizontal = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  sprite58ScaleUpVertical = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  sprite59ScaleUpHorizontal = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  sprite59ScaleUpVertical = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  sprite60ScaleUpHorizontal = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  sprite60ScaleUpVertical = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  viewBoxXReg = _RAND_193[9:0];
  _RAND_194 = {1{`RANDOM}};
  viewBoxYReg = _RAND_194[8:0];
  _RAND_195 = {1{`RANDOM}};
  lvlReg = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  livesReg = _RAND_196[2:0];
  _RAND_197 = {1{`RANDOM}};
  extraLifeCnt = _RAND_197[9:0];
  _RAND_198 = {1{`RANDOM}};
  spawnDelayCounter = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  nextSpriteToSpawn = _RAND_199[5:0];
  _RAND_200 = {1{`RANDOM}};
  starCnt = _RAND_200[9:0];
  _RAND_201 = {1{`RANDOM}};
  collisionDetected = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  blinkCounter = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  blinkTimes = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  isBlinking = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  spriteXRegs_58_REG = _RAND_205[10:0];
  _RAND_206 = {1{`RANDOM}};
  spriteYRegs_58_REG = _RAND_206[9:0];
  _RAND_207 = {1{`RANDOM}};
  spriteXRegs_59_REG = _RAND_207[10:0];
  _RAND_208 = {1{`RANDOM}};
  spriteYRegs_59_REG = _RAND_208[9:0];
  _RAND_209 = {1{`RANDOM}};
  spriteXRegs_60_REG = _RAND_209[10:0];
  _RAND_210 = {1{`RANDOM}};
  spriteYRegs_60_REG = _RAND_210[9:0];
  _RAND_211 = {1{`RANDOM}};
  spriteXRegs_58_REG_1 = _RAND_211[10:0];
  _RAND_212 = {1{`RANDOM}};
  spriteYRegs_58_REG_1 = _RAND_212[9:0];
  _RAND_213 = {1{`RANDOM}};
  spriteXRegs_59_REG_1 = _RAND_213[10:0];
  _RAND_214 = {1{`RANDOM}};
  spriteYRegs_59_REG_1 = _RAND_214[9:0];
  _RAND_215 = {1{`RANDOM}};
  spriteXRegs_60_REG_1 = _RAND_215[10:0];
  _RAND_216 = {1{`RANDOM}};
  spriteYRegs_60_REG_1 = _RAND_216[9:0];
  _RAND_217 = {1{`RANDOM}};
  spriteXRegs_58_REG_2 = _RAND_217[10:0];
  _RAND_218 = {1{`RANDOM}};
  spriteYRegs_58_REG_2 = _RAND_218[9:0];
  _RAND_219 = {1{`RANDOM}};
  spriteXRegs_59_REG_2 = _RAND_219[10:0];
  _RAND_220 = {1{`RANDOM}};
  spriteYRegs_59_REG_2 = _RAND_220[9:0];
  _RAND_221 = {1{`RANDOM}};
  spriteXRegs_60_REG_2 = _RAND_221[10:0];
  _RAND_222 = {1{`RANDOM}};
  spriteYRegs_60_REG_2 = _RAND_222[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GameTop(
  input        clock,
  input        reset,
  input        io_btnC, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnU, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnL, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnR, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnD, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaRed, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaBlue, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaGreen, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_Hsync, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_Vsync, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_missingFrameError, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_viewBoxOutOfRangeError // @[\\src\\main\\scala\\GameTop.scala 14:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  graphicEngineVGA_clock; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_reset; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_46; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_47; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_48; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_49; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_50; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_51; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_52; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_53; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_54; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_55; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_56; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_57; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_61; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_62; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_63; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_46; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_47; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_48; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_49; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_50; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_51; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_52; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_53; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_54; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_55; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_56; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_57; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_61; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_62; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_63; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_46; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_47; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_48; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_49; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_50; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_51; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_52; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_53; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_54; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_55; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_56; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_57; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_61; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_62; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_63; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [8:0] graphicEngineVGA_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_missingFrameError; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaRed; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaBlue; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaGreen; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Hsync; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Vsync; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  soundEngine_clock; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  soundEngine_reset; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  gameLogic_clock; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_reset; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnC; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnU; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnL; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnR; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnD; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_46; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_47; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_48; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_49; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_50; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_51; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_52; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_53; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_54; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_55; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_56; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_57; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_61; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_62; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_63; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_46; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_47; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_48; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_49; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_50; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_51; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_52; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_53; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_54; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_55; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_56; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_57; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_61; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_62; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_63; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_46; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_47; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_48; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_49; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_50; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_51; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_52; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_53; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_54; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_55; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_56; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_57; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_61; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_62; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_63; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [8:0] gameLogic_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  reg [20:0] debounceCounter; // @[\\src\\main\\scala\\GameTop.scala 68:32]
  wire  debounceSampleEn = debounceCounter == 21'h1e847f; // @[\\src\\main\\scala\\GameTop.scala 70:24]
  wire [20:0] _debounceCounter_T_1 = debounceCounter + 21'h1; // @[\\src\\main\\scala\\GameTop.scala 74:40]
  reg [21:0] resetReleaseCounter; // @[\\src\\main\\scala\\GameTop.scala 81:36]
  wire [21:0] _resetReleaseCounter_T_1 = resetReleaseCounter + 22'h1; // @[\\src\\main\\scala\\GameTop.scala 87:48]
  reg  btnCState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnCState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnCState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnCState; // @[\\src\\main\\scala\\GameTop.scala 93:28]
  reg  btnUState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState; // @[\\src\\main\\scala\\GameTop.scala 94:28]
  reg  btnLState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState; // @[\\src\\main\\scala\\GameTop.scala 95:28]
  reg  btnRState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState; // @[\\src\\main\\scala\\GameTop.scala 96:28]
  reg  btnDState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState; // @[\\src\\main\\scala\\GameTop.scala 97:28]
  GraphicEngineVGA graphicEngineVGA ( // @[\\src\\main\\scala\\GameTop.scala 46:32]
    .clock(graphicEngineVGA_clock),
    .reset(graphicEngineVGA_reset),
    .io_spriteXPosition_3(graphicEngineVGA_io_spriteXPosition_3),
    .io_spriteXPosition_7(graphicEngineVGA_io_spriteXPosition_7),
    .io_spriteXPosition_8(graphicEngineVGA_io_spriteXPosition_8),
    .io_spriteXPosition_9(graphicEngineVGA_io_spriteXPosition_9),
    .io_spriteXPosition_10(graphicEngineVGA_io_spriteXPosition_10),
    .io_spriteXPosition_11(graphicEngineVGA_io_spriteXPosition_11),
    .io_spriteXPosition_12(graphicEngineVGA_io_spriteXPosition_12),
    .io_spriteXPosition_13(graphicEngineVGA_io_spriteXPosition_13),
    .io_spriteXPosition_14(graphicEngineVGA_io_spriteXPosition_14),
    .io_spriteXPosition_16(graphicEngineVGA_io_spriteXPosition_16),
    .io_spriteXPosition_17(graphicEngineVGA_io_spriteXPosition_17),
    .io_spriteXPosition_18(graphicEngineVGA_io_spriteXPosition_18),
    .io_spriteXPosition_19(graphicEngineVGA_io_spriteXPosition_19),
    .io_spriteXPosition_20(graphicEngineVGA_io_spriteXPosition_20),
    .io_spriteXPosition_21(graphicEngineVGA_io_spriteXPosition_21),
    .io_spriteXPosition_22(graphicEngineVGA_io_spriteXPosition_22),
    .io_spriteXPosition_23(graphicEngineVGA_io_spriteXPosition_23),
    .io_spriteXPosition_24(graphicEngineVGA_io_spriteXPosition_24),
    .io_spriteXPosition_25(graphicEngineVGA_io_spriteXPosition_25),
    .io_spriteXPosition_26(graphicEngineVGA_io_spriteXPosition_26),
    .io_spriteXPosition_27(graphicEngineVGA_io_spriteXPosition_27),
    .io_spriteXPosition_28(graphicEngineVGA_io_spriteXPosition_28),
    .io_spriteXPosition_29(graphicEngineVGA_io_spriteXPosition_29),
    .io_spriteXPosition_30(graphicEngineVGA_io_spriteXPosition_30),
    .io_spriteXPosition_31(graphicEngineVGA_io_spriteXPosition_31),
    .io_spriteXPosition_32(graphicEngineVGA_io_spriteXPosition_32),
    .io_spriteXPosition_33(graphicEngineVGA_io_spriteXPosition_33),
    .io_spriteXPosition_34(graphicEngineVGA_io_spriteXPosition_34),
    .io_spriteXPosition_35(graphicEngineVGA_io_spriteXPosition_35),
    .io_spriteXPosition_36(graphicEngineVGA_io_spriteXPosition_36),
    .io_spriteXPosition_37(graphicEngineVGA_io_spriteXPosition_37),
    .io_spriteXPosition_38(graphicEngineVGA_io_spriteXPosition_38),
    .io_spriteXPosition_39(graphicEngineVGA_io_spriteXPosition_39),
    .io_spriteXPosition_40(graphicEngineVGA_io_spriteXPosition_40),
    .io_spriteXPosition_41(graphicEngineVGA_io_spriteXPosition_41),
    .io_spriteXPosition_42(graphicEngineVGA_io_spriteXPosition_42),
    .io_spriteXPosition_43(graphicEngineVGA_io_spriteXPosition_43),
    .io_spriteXPosition_44(graphicEngineVGA_io_spriteXPosition_44),
    .io_spriteXPosition_45(graphicEngineVGA_io_spriteXPosition_45),
    .io_spriteXPosition_46(graphicEngineVGA_io_spriteXPosition_46),
    .io_spriteXPosition_47(graphicEngineVGA_io_spriteXPosition_47),
    .io_spriteXPosition_48(graphicEngineVGA_io_spriteXPosition_48),
    .io_spriteXPosition_49(graphicEngineVGA_io_spriteXPosition_49),
    .io_spriteXPosition_50(graphicEngineVGA_io_spriteXPosition_50),
    .io_spriteXPosition_51(graphicEngineVGA_io_spriteXPosition_51),
    .io_spriteXPosition_52(graphicEngineVGA_io_spriteXPosition_52),
    .io_spriteXPosition_53(graphicEngineVGA_io_spriteXPosition_53),
    .io_spriteXPosition_54(graphicEngineVGA_io_spriteXPosition_54),
    .io_spriteXPosition_55(graphicEngineVGA_io_spriteXPosition_55),
    .io_spriteXPosition_56(graphicEngineVGA_io_spriteXPosition_56),
    .io_spriteXPosition_57(graphicEngineVGA_io_spriteXPosition_57),
    .io_spriteXPosition_58(graphicEngineVGA_io_spriteXPosition_58),
    .io_spriteXPosition_59(graphicEngineVGA_io_spriteXPosition_59),
    .io_spriteXPosition_60(graphicEngineVGA_io_spriteXPosition_60),
    .io_spriteXPosition_61(graphicEngineVGA_io_spriteXPosition_61),
    .io_spriteXPosition_62(graphicEngineVGA_io_spriteXPosition_62),
    .io_spriteXPosition_63(graphicEngineVGA_io_spriteXPosition_63),
    .io_spriteYPosition_3(graphicEngineVGA_io_spriteYPosition_3),
    .io_spriteYPosition_7(graphicEngineVGA_io_spriteYPosition_7),
    .io_spriteYPosition_8(graphicEngineVGA_io_spriteYPosition_8),
    .io_spriteYPosition_9(graphicEngineVGA_io_spriteYPosition_9),
    .io_spriteYPosition_10(graphicEngineVGA_io_spriteYPosition_10),
    .io_spriteYPosition_11(graphicEngineVGA_io_spriteYPosition_11),
    .io_spriteYPosition_12(graphicEngineVGA_io_spriteYPosition_12),
    .io_spriteYPosition_13(graphicEngineVGA_io_spriteYPosition_13),
    .io_spriteYPosition_14(graphicEngineVGA_io_spriteYPosition_14),
    .io_spriteYPosition_16(graphicEngineVGA_io_spriteYPosition_16),
    .io_spriteYPosition_17(graphicEngineVGA_io_spriteYPosition_17),
    .io_spriteYPosition_18(graphicEngineVGA_io_spriteYPosition_18),
    .io_spriteYPosition_19(graphicEngineVGA_io_spriteYPosition_19),
    .io_spriteYPosition_20(graphicEngineVGA_io_spriteYPosition_20),
    .io_spriteYPosition_21(graphicEngineVGA_io_spriteYPosition_21),
    .io_spriteYPosition_22(graphicEngineVGA_io_spriteYPosition_22),
    .io_spriteYPosition_23(graphicEngineVGA_io_spriteYPosition_23),
    .io_spriteYPosition_24(graphicEngineVGA_io_spriteYPosition_24),
    .io_spriteYPosition_25(graphicEngineVGA_io_spriteYPosition_25),
    .io_spriteYPosition_26(graphicEngineVGA_io_spriteYPosition_26),
    .io_spriteYPosition_27(graphicEngineVGA_io_spriteYPosition_27),
    .io_spriteYPosition_28(graphicEngineVGA_io_spriteYPosition_28),
    .io_spriteYPosition_29(graphicEngineVGA_io_spriteYPosition_29),
    .io_spriteYPosition_30(graphicEngineVGA_io_spriteYPosition_30),
    .io_spriteYPosition_31(graphicEngineVGA_io_spriteYPosition_31),
    .io_spriteYPosition_32(graphicEngineVGA_io_spriteYPosition_32),
    .io_spriteYPosition_33(graphicEngineVGA_io_spriteYPosition_33),
    .io_spriteYPosition_34(graphicEngineVGA_io_spriteYPosition_34),
    .io_spriteYPosition_35(graphicEngineVGA_io_spriteYPosition_35),
    .io_spriteYPosition_36(graphicEngineVGA_io_spriteYPosition_36),
    .io_spriteYPosition_37(graphicEngineVGA_io_spriteYPosition_37),
    .io_spriteYPosition_38(graphicEngineVGA_io_spriteYPosition_38),
    .io_spriteYPosition_39(graphicEngineVGA_io_spriteYPosition_39),
    .io_spriteYPosition_40(graphicEngineVGA_io_spriteYPosition_40),
    .io_spriteYPosition_41(graphicEngineVGA_io_spriteYPosition_41),
    .io_spriteYPosition_42(graphicEngineVGA_io_spriteYPosition_42),
    .io_spriteYPosition_43(graphicEngineVGA_io_spriteYPosition_43),
    .io_spriteYPosition_44(graphicEngineVGA_io_spriteYPosition_44),
    .io_spriteYPosition_45(graphicEngineVGA_io_spriteYPosition_45),
    .io_spriteYPosition_46(graphicEngineVGA_io_spriteYPosition_46),
    .io_spriteYPosition_47(graphicEngineVGA_io_spriteYPosition_47),
    .io_spriteYPosition_48(graphicEngineVGA_io_spriteYPosition_48),
    .io_spriteYPosition_49(graphicEngineVGA_io_spriteYPosition_49),
    .io_spriteYPosition_50(graphicEngineVGA_io_spriteYPosition_50),
    .io_spriteYPosition_51(graphicEngineVGA_io_spriteYPosition_51),
    .io_spriteYPosition_52(graphicEngineVGA_io_spriteYPosition_52),
    .io_spriteYPosition_53(graphicEngineVGA_io_spriteYPosition_53),
    .io_spriteYPosition_54(graphicEngineVGA_io_spriteYPosition_54),
    .io_spriteYPosition_55(graphicEngineVGA_io_spriteYPosition_55),
    .io_spriteYPosition_56(graphicEngineVGA_io_spriteYPosition_56),
    .io_spriteYPosition_57(graphicEngineVGA_io_spriteYPosition_57),
    .io_spriteYPosition_58(graphicEngineVGA_io_spriteYPosition_58),
    .io_spriteYPosition_59(graphicEngineVGA_io_spriteYPosition_59),
    .io_spriteYPosition_60(graphicEngineVGA_io_spriteYPosition_60),
    .io_spriteYPosition_61(graphicEngineVGA_io_spriteYPosition_61),
    .io_spriteYPosition_62(graphicEngineVGA_io_spriteYPosition_62),
    .io_spriteYPosition_63(graphicEngineVGA_io_spriteYPosition_63),
    .io_spriteVisible_3(graphicEngineVGA_io_spriteVisible_3),
    .io_spriteVisible_4(graphicEngineVGA_io_spriteVisible_4),
    .io_spriteVisible_5(graphicEngineVGA_io_spriteVisible_5),
    .io_spriteVisible_6(graphicEngineVGA_io_spriteVisible_6),
    .io_spriteVisible_7(graphicEngineVGA_io_spriteVisible_7),
    .io_spriteVisible_8(graphicEngineVGA_io_spriteVisible_8),
    .io_spriteVisible_9(graphicEngineVGA_io_spriteVisible_9),
    .io_spriteVisible_10(graphicEngineVGA_io_spriteVisible_10),
    .io_spriteVisible_11(graphicEngineVGA_io_spriteVisible_11),
    .io_spriteVisible_12(graphicEngineVGA_io_spriteVisible_12),
    .io_spriteVisible_13(graphicEngineVGA_io_spriteVisible_13),
    .io_spriteVisible_14(graphicEngineVGA_io_spriteVisible_14),
    .io_spriteVisible_15(graphicEngineVGA_io_spriteVisible_15),
    .io_spriteVisible_16(graphicEngineVGA_io_spriteVisible_16),
    .io_spriteVisible_17(graphicEngineVGA_io_spriteVisible_17),
    .io_spriteVisible_18(graphicEngineVGA_io_spriteVisible_18),
    .io_spriteVisible_19(graphicEngineVGA_io_spriteVisible_19),
    .io_spriteVisible_20(graphicEngineVGA_io_spriteVisible_20),
    .io_spriteVisible_21(graphicEngineVGA_io_spriteVisible_21),
    .io_spriteVisible_22(graphicEngineVGA_io_spriteVisible_22),
    .io_spriteVisible_23(graphicEngineVGA_io_spriteVisible_23),
    .io_spriteVisible_24(graphicEngineVGA_io_spriteVisible_24),
    .io_spriteVisible_25(graphicEngineVGA_io_spriteVisible_25),
    .io_spriteVisible_26(graphicEngineVGA_io_spriteVisible_26),
    .io_spriteVisible_27(graphicEngineVGA_io_spriteVisible_27),
    .io_spriteVisible_28(graphicEngineVGA_io_spriteVisible_28),
    .io_spriteVisible_29(graphicEngineVGA_io_spriteVisible_29),
    .io_spriteVisible_30(graphicEngineVGA_io_spriteVisible_30),
    .io_spriteVisible_31(graphicEngineVGA_io_spriteVisible_31),
    .io_spriteVisible_32(graphicEngineVGA_io_spriteVisible_32),
    .io_spriteVisible_33(graphicEngineVGA_io_spriteVisible_33),
    .io_spriteVisible_34(graphicEngineVGA_io_spriteVisible_34),
    .io_spriteVisible_35(graphicEngineVGA_io_spriteVisible_35),
    .io_spriteVisible_36(graphicEngineVGA_io_spriteVisible_36),
    .io_spriteVisible_37(graphicEngineVGA_io_spriteVisible_37),
    .io_spriteVisible_38(graphicEngineVGA_io_spriteVisible_38),
    .io_spriteVisible_39(graphicEngineVGA_io_spriteVisible_39),
    .io_spriteVisible_40(graphicEngineVGA_io_spriteVisible_40),
    .io_spriteVisible_41(graphicEngineVGA_io_spriteVisible_41),
    .io_spriteVisible_42(graphicEngineVGA_io_spriteVisible_42),
    .io_spriteVisible_43(graphicEngineVGA_io_spriteVisible_43),
    .io_spriteVisible_44(graphicEngineVGA_io_spriteVisible_44),
    .io_spriteVisible_45(graphicEngineVGA_io_spriteVisible_45),
    .io_spriteVisible_46(graphicEngineVGA_io_spriteVisible_46),
    .io_spriteVisible_47(graphicEngineVGA_io_spriteVisible_47),
    .io_spriteVisible_48(graphicEngineVGA_io_spriteVisible_48),
    .io_spriteVisible_49(graphicEngineVGA_io_spriteVisible_49),
    .io_spriteVisible_50(graphicEngineVGA_io_spriteVisible_50),
    .io_spriteVisible_51(graphicEngineVGA_io_spriteVisible_51),
    .io_spriteVisible_52(graphicEngineVGA_io_spriteVisible_52),
    .io_spriteVisible_53(graphicEngineVGA_io_spriteVisible_53),
    .io_spriteVisible_54(graphicEngineVGA_io_spriteVisible_54),
    .io_spriteVisible_55(graphicEngineVGA_io_spriteVisible_55),
    .io_spriteVisible_56(graphicEngineVGA_io_spriteVisible_56),
    .io_spriteVisible_57(graphicEngineVGA_io_spriteVisible_57),
    .io_spriteVisible_58(graphicEngineVGA_io_spriteVisible_58),
    .io_spriteVisible_59(graphicEngineVGA_io_spriteVisible_59),
    .io_spriteVisible_60(graphicEngineVGA_io_spriteVisible_60),
    .io_spriteVisible_61(graphicEngineVGA_io_spriteVisible_61),
    .io_spriteVisible_62(graphicEngineVGA_io_spriteVisible_62),
    .io_spriteVisible_63(graphicEngineVGA_io_spriteVisible_63),
    .io_spriteScaleUpHorizontal_16(graphicEngineVGA_io_spriteScaleUpHorizontal_16),
    .io_spriteScaleUpHorizontal_17(graphicEngineVGA_io_spriteScaleUpHorizontal_17),
    .io_spriteScaleUpHorizontal_18(graphicEngineVGA_io_spriteScaleUpHorizontal_18),
    .io_spriteScaleUpHorizontal_19(graphicEngineVGA_io_spriteScaleUpHorizontal_19),
    .io_spriteScaleUpHorizontal_20(graphicEngineVGA_io_spriteScaleUpHorizontal_20),
    .io_spriteScaleUpHorizontal_21(graphicEngineVGA_io_spriteScaleUpHorizontal_21),
    .io_spriteScaleUpHorizontal_22(graphicEngineVGA_io_spriteScaleUpHorizontal_22),
    .io_spriteScaleUpHorizontal_23(graphicEngineVGA_io_spriteScaleUpHorizontal_23),
    .io_spriteScaleUpHorizontal_24(graphicEngineVGA_io_spriteScaleUpHorizontal_24),
    .io_spriteScaleUpHorizontal_25(graphicEngineVGA_io_spriteScaleUpHorizontal_25),
    .io_spriteScaleUpHorizontal_26(graphicEngineVGA_io_spriteScaleUpHorizontal_26),
    .io_spriteScaleUpHorizontal_27(graphicEngineVGA_io_spriteScaleUpHorizontal_27),
    .io_spriteScaleUpHorizontal_28(graphicEngineVGA_io_spriteScaleUpHorizontal_28),
    .io_spriteScaleUpHorizontal_29(graphicEngineVGA_io_spriteScaleUpHorizontal_29),
    .io_spriteScaleUpHorizontal_30(graphicEngineVGA_io_spriteScaleUpHorizontal_30),
    .io_spriteScaleUpHorizontal_31(graphicEngineVGA_io_spriteScaleUpHorizontal_31),
    .io_spriteScaleUpHorizontal_32(graphicEngineVGA_io_spriteScaleUpHorizontal_32),
    .io_spriteScaleUpHorizontal_33(graphicEngineVGA_io_spriteScaleUpHorizontal_33),
    .io_spriteScaleUpHorizontal_34(graphicEngineVGA_io_spriteScaleUpHorizontal_34),
    .io_spriteScaleUpHorizontal_35(graphicEngineVGA_io_spriteScaleUpHorizontal_35),
    .io_spriteScaleUpHorizontal_36(graphicEngineVGA_io_spriteScaleUpHorizontal_36),
    .io_spriteScaleUpHorizontal_37(graphicEngineVGA_io_spriteScaleUpHorizontal_37),
    .io_spriteScaleUpHorizontal_38(graphicEngineVGA_io_spriteScaleUpHorizontal_38),
    .io_spriteScaleUpHorizontal_39(graphicEngineVGA_io_spriteScaleUpHorizontal_39),
    .io_spriteScaleUpHorizontal_40(graphicEngineVGA_io_spriteScaleUpHorizontal_40),
    .io_spriteScaleUpHorizontal_41(graphicEngineVGA_io_spriteScaleUpHorizontal_41),
    .io_spriteScaleUpHorizontal_42(graphicEngineVGA_io_spriteScaleUpHorizontal_42),
    .io_spriteScaleUpHorizontal_43(graphicEngineVGA_io_spriteScaleUpHorizontal_43),
    .io_spriteScaleUpHorizontal_44(graphicEngineVGA_io_spriteScaleUpHorizontal_44),
    .io_spriteScaleUpHorizontal_45(graphicEngineVGA_io_spriteScaleUpHorizontal_45),
    .io_spriteScaleUpHorizontal_58(graphicEngineVGA_io_spriteScaleUpHorizontal_58),
    .io_spriteScaleUpHorizontal_59(graphicEngineVGA_io_spriteScaleUpHorizontal_59),
    .io_spriteScaleUpHorizontal_60(graphicEngineVGA_io_spriteScaleUpHorizontal_60),
    .io_spriteScaleUpVertical_16(graphicEngineVGA_io_spriteScaleUpVertical_16),
    .io_spriteScaleUpVertical_17(graphicEngineVGA_io_spriteScaleUpVertical_17),
    .io_spriteScaleUpVertical_18(graphicEngineVGA_io_spriteScaleUpVertical_18),
    .io_spriteScaleUpVertical_19(graphicEngineVGA_io_spriteScaleUpVertical_19),
    .io_spriteScaleUpVertical_20(graphicEngineVGA_io_spriteScaleUpVertical_20),
    .io_spriteScaleUpVertical_21(graphicEngineVGA_io_spriteScaleUpVertical_21),
    .io_spriteScaleUpVertical_22(graphicEngineVGA_io_spriteScaleUpVertical_22),
    .io_spriteScaleUpVertical_23(graphicEngineVGA_io_spriteScaleUpVertical_23),
    .io_spriteScaleUpVertical_24(graphicEngineVGA_io_spriteScaleUpVertical_24),
    .io_spriteScaleUpVertical_25(graphicEngineVGA_io_spriteScaleUpVertical_25),
    .io_spriteScaleUpVertical_26(graphicEngineVGA_io_spriteScaleUpVertical_26),
    .io_spriteScaleUpVertical_27(graphicEngineVGA_io_spriteScaleUpVertical_27),
    .io_spriteScaleUpVertical_28(graphicEngineVGA_io_spriteScaleUpVertical_28),
    .io_spriteScaleUpVertical_29(graphicEngineVGA_io_spriteScaleUpVertical_29),
    .io_spriteScaleUpVertical_30(graphicEngineVGA_io_spriteScaleUpVertical_30),
    .io_spriteScaleUpVertical_31(graphicEngineVGA_io_spriteScaleUpVertical_31),
    .io_spriteScaleUpVertical_32(graphicEngineVGA_io_spriteScaleUpVertical_32),
    .io_spriteScaleUpVertical_33(graphicEngineVGA_io_spriteScaleUpVertical_33),
    .io_spriteScaleUpVertical_34(graphicEngineVGA_io_spriteScaleUpVertical_34),
    .io_spriteScaleUpVertical_35(graphicEngineVGA_io_spriteScaleUpVertical_35),
    .io_spriteScaleUpVertical_36(graphicEngineVGA_io_spriteScaleUpVertical_36),
    .io_spriteScaleUpVertical_37(graphicEngineVGA_io_spriteScaleUpVertical_37),
    .io_spriteScaleUpVertical_38(graphicEngineVGA_io_spriteScaleUpVertical_38),
    .io_spriteScaleUpVertical_39(graphicEngineVGA_io_spriteScaleUpVertical_39),
    .io_spriteScaleUpVertical_40(graphicEngineVGA_io_spriteScaleUpVertical_40),
    .io_spriteScaleUpVertical_41(graphicEngineVGA_io_spriteScaleUpVertical_41),
    .io_spriteScaleUpVertical_42(graphicEngineVGA_io_spriteScaleUpVertical_42),
    .io_spriteScaleUpVertical_43(graphicEngineVGA_io_spriteScaleUpVertical_43),
    .io_spriteScaleUpVertical_44(graphicEngineVGA_io_spriteScaleUpVertical_44),
    .io_spriteScaleUpVertical_45(graphicEngineVGA_io_spriteScaleUpVertical_45),
    .io_spriteScaleUpVertical_58(graphicEngineVGA_io_spriteScaleUpVertical_58),
    .io_spriteScaleUpVertical_59(graphicEngineVGA_io_spriteScaleUpVertical_59),
    .io_spriteScaleUpVertical_60(graphicEngineVGA_io_spriteScaleUpVertical_60),
    .io_viewBoxX(graphicEngineVGA_io_viewBoxX),
    .io_viewBoxY(graphicEngineVGA_io_viewBoxY),
    .io_newFrame(graphicEngineVGA_io_newFrame),
    .io_frameUpdateDone(graphicEngineVGA_io_frameUpdateDone),
    .io_missingFrameError(graphicEngineVGA_io_missingFrameError),
    .io_viewBoxOutOfRangeError(graphicEngineVGA_io_viewBoxOutOfRangeError),
    .io_vgaRed(graphicEngineVGA_io_vgaRed),
    .io_vgaBlue(graphicEngineVGA_io_vgaBlue),
    .io_vgaGreen(graphicEngineVGA_io_vgaGreen),
    .io_Hsync(graphicEngineVGA_io_Hsync),
    .io_Vsync(graphicEngineVGA_io_Vsync)
  );
  SoundEngine soundEngine ( // @[\\src\\main\\scala\\GameTop.scala 49:27]
    .clock(soundEngine_clock),
    .reset(soundEngine_reset)
  );
  GameLogic gameLogic ( // @[\\src\\main\\scala\\GameTop.scala 53:25]
    .clock(gameLogic_clock),
    .reset(gameLogic_reset),
    .io_btnC(gameLogic_io_btnC),
    .io_btnU(gameLogic_io_btnU),
    .io_btnL(gameLogic_io_btnL),
    .io_btnR(gameLogic_io_btnR),
    .io_btnD(gameLogic_io_btnD),
    .io_spriteXPosition_3(gameLogic_io_spriteXPosition_3),
    .io_spriteXPosition_7(gameLogic_io_spriteXPosition_7),
    .io_spriteXPosition_8(gameLogic_io_spriteXPosition_8),
    .io_spriteXPosition_9(gameLogic_io_spriteXPosition_9),
    .io_spriteXPosition_10(gameLogic_io_spriteXPosition_10),
    .io_spriteXPosition_11(gameLogic_io_spriteXPosition_11),
    .io_spriteXPosition_12(gameLogic_io_spriteXPosition_12),
    .io_spriteXPosition_13(gameLogic_io_spriteXPosition_13),
    .io_spriteXPosition_14(gameLogic_io_spriteXPosition_14),
    .io_spriteXPosition_16(gameLogic_io_spriteXPosition_16),
    .io_spriteXPosition_17(gameLogic_io_spriteXPosition_17),
    .io_spriteXPosition_18(gameLogic_io_spriteXPosition_18),
    .io_spriteXPosition_19(gameLogic_io_spriteXPosition_19),
    .io_spriteXPosition_20(gameLogic_io_spriteXPosition_20),
    .io_spriteXPosition_21(gameLogic_io_spriteXPosition_21),
    .io_spriteXPosition_22(gameLogic_io_spriteXPosition_22),
    .io_spriteXPosition_23(gameLogic_io_spriteXPosition_23),
    .io_spriteXPosition_24(gameLogic_io_spriteXPosition_24),
    .io_spriteXPosition_25(gameLogic_io_spriteXPosition_25),
    .io_spriteXPosition_26(gameLogic_io_spriteXPosition_26),
    .io_spriteXPosition_27(gameLogic_io_spriteXPosition_27),
    .io_spriteXPosition_28(gameLogic_io_spriteXPosition_28),
    .io_spriteXPosition_29(gameLogic_io_spriteXPosition_29),
    .io_spriteXPosition_30(gameLogic_io_spriteXPosition_30),
    .io_spriteXPosition_31(gameLogic_io_spriteXPosition_31),
    .io_spriteXPosition_32(gameLogic_io_spriteXPosition_32),
    .io_spriteXPosition_33(gameLogic_io_spriteXPosition_33),
    .io_spriteXPosition_34(gameLogic_io_spriteXPosition_34),
    .io_spriteXPosition_35(gameLogic_io_spriteXPosition_35),
    .io_spriteXPosition_36(gameLogic_io_spriteXPosition_36),
    .io_spriteXPosition_37(gameLogic_io_spriteXPosition_37),
    .io_spriteXPosition_38(gameLogic_io_spriteXPosition_38),
    .io_spriteXPosition_39(gameLogic_io_spriteXPosition_39),
    .io_spriteXPosition_40(gameLogic_io_spriteXPosition_40),
    .io_spriteXPosition_41(gameLogic_io_spriteXPosition_41),
    .io_spriteXPosition_42(gameLogic_io_spriteXPosition_42),
    .io_spriteXPosition_43(gameLogic_io_spriteXPosition_43),
    .io_spriteXPosition_44(gameLogic_io_spriteXPosition_44),
    .io_spriteXPosition_45(gameLogic_io_spriteXPosition_45),
    .io_spriteXPosition_46(gameLogic_io_spriteXPosition_46),
    .io_spriteXPosition_47(gameLogic_io_spriteXPosition_47),
    .io_spriteXPosition_48(gameLogic_io_spriteXPosition_48),
    .io_spriteXPosition_49(gameLogic_io_spriteXPosition_49),
    .io_spriteXPosition_50(gameLogic_io_spriteXPosition_50),
    .io_spriteXPosition_51(gameLogic_io_spriteXPosition_51),
    .io_spriteXPosition_52(gameLogic_io_spriteXPosition_52),
    .io_spriteXPosition_53(gameLogic_io_spriteXPosition_53),
    .io_spriteXPosition_54(gameLogic_io_spriteXPosition_54),
    .io_spriteXPosition_55(gameLogic_io_spriteXPosition_55),
    .io_spriteXPosition_56(gameLogic_io_spriteXPosition_56),
    .io_spriteXPosition_57(gameLogic_io_spriteXPosition_57),
    .io_spriteXPosition_58(gameLogic_io_spriteXPosition_58),
    .io_spriteXPosition_59(gameLogic_io_spriteXPosition_59),
    .io_spriteXPosition_60(gameLogic_io_spriteXPosition_60),
    .io_spriteXPosition_61(gameLogic_io_spriteXPosition_61),
    .io_spriteXPosition_62(gameLogic_io_spriteXPosition_62),
    .io_spriteXPosition_63(gameLogic_io_spriteXPosition_63),
    .io_spriteYPosition_3(gameLogic_io_spriteYPosition_3),
    .io_spriteYPosition_7(gameLogic_io_spriteYPosition_7),
    .io_spriteYPosition_8(gameLogic_io_spriteYPosition_8),
    .io_spriteYPosition_9(gameLogic_io_spriteYPosition_9),
    .io_spriteYPosition_10(gameLogic_io_spriteYPosition_10),
    .io_spriteYPosition_11(gameLogic_io_spriteYPosition_11),
    .io_spriteYPosition_12(gameLogic_io_spriteYPosition_12),
    .io_spriteYPosition_13(gameLogic_io_spriteYPosition_13),
    .io_spriteYPosition_14(gameLogic_io_spriteYPosition_14),
    .io_spriteYPosition_16(gameLogic_io_spriteYPosition_16),
    .io_spriteYPosition_17(gameLogic_io_spriteYPosition_17),
    .io_spriteYPosition_18(gameLogic_io_spriteYPosition_18),
    .io_spriteYPosition_19(gameLogic_io_spriteYPosition_19),
    .io_spriteYPosition_20(gameLogic_io_spriteYPosition_20),
    .io_spriteYPosition_21(gameLogic_io_spriteYPosition_21),
    .io_spriteYPosition_22(gameLogic_io_spriteYPosition_22),
    .io_spriteYPosition_23(gameLogic_io_spriteYPosition_23),
    .io_spriteYPosition_24(gameLogic_io_spriteYPosition_24),
    .io_spriteYPosition_25(gameLogic_io_spriteYPosition_25),
    .io_spriteYPosition_26(gameLogic_io_spriteYPosition_26),
    .io_spriteYPosition_27(gameLogic_io_spriteYPosition_27),
    .io_spriteYPosition_28(gameLogic_io_spriteYPosition_28),
    .io_spriteYPosition_29(gameLogic_io_spriteYPosition_29),
    .io_spriteYPosition_30(gameLogic_io_spriteYPosition_30),
    .io_spriteYPosition_31(gameLogic_io_spriteYPosition_31),
    .io_spriteYPosition_32(gameLogic_io_spriteYPosition_32),
    .io_spriteYPosition_33(gameLogic_io_spriteYPosition_33),
    .io_spriteYPosition_34(gameLogic_io_spriteYPosition_34),
    .io_spriteYPosition_35(gameLogic_io_spriteYPosition_35),
    .io_spriteYPosition_36(gameLogic_io_spriteYPosition_36),
    .io_spriteYPosition_37(gameLogic_io_spriteYPosition_37),
    .io_spriteYPosition_38(gameLogic_io_spriteYPosition_38),
    .io_spriteYPosition_39(gameLogic_io_spriteYPosition_39),
    .io_spriteYPosition_40(gameLogic_io_spriteYPosition_40),
    .io_spriteYPosition_41(gameLogic_io_spriteYPosition_41),
    .io_spriteYPosition_42(gameLogic_io_spriteYPosition_42),
    .io_spriteYPosition_43(gameLogic_io_spriteYPosition_43),
    .io_spriteYPosition_44(gameLogic_io_spriteYPosition_44),
    .io_spriteYPosition_45(gameLogic_io_spriteYPosition_45),
    .io_spriteYPosition_46(gameLogic_io_spriteYPosition_46),
    .io_spriteYPosition_47(gameLogic_io_spriteYPosition_47),
    .io_spriteYPosition_48(gameLogic_io_spriteYPosition_48),
    .io_spriteYPosition_49(gameLogic_io_spriteYPosition_49),
    .io_spriteYPosition_50(gameLogic_io_spriteYPosition_50),
    .io_spriteYPosition_51(gameLogic_io_spriteYPosition_51),
    .io_spriteYPosition_52(gameLogic_io_spriteYPosition_52),
    .io_spriteYPosition_53(gameLogic_io_spriteYPosition_53),
    .io_spriteYPosition_54(gameLogic_io_spriteYPosition_54),
    .io_spriteYPosition_55(gameLogic_io_spriteYPosition_55),
    .io_spriteYPosition_56(gameLogic_io_spriteYPosition_56),
    .io_spriteYPosition_57(gameLogic_io_spriteYPosition_57),
    .io_spriteYPosition_58(gameLogic_io_spriteYPosition_58),
    .io_spriteYPosition_59(gameLogic_io_spriteYPosition_59),
    .io_spriteYPosition_60(gameLogic_io_spriteYPosition_60),
    .io_spriteYPosition_61(gameLogic_io_spriteYPosition_61),
    .io_spriteYPosition_62(gameLogic_io_spriteYPosition_62),
    .io_spriteYPosition_63(gameLogic_io_spriteYPosition_63),
    .io_spriteVisible_3(gameLogic_io_spriteVisible_3),
    .io_spriteVisible_4(gameLogic_io_spriteVisible_4),
    .io_spriteVisible_5(gameLogic_io_spriteVisible_5),
    .io_spriteVisible_6(gameLogic_io_spriteVisible_6),
    .io_spriteVisible_7(gameLogic_io_spriteVisible_7),
    .io_spriteVisible_8(gameLogic_io_spriteVisible_8),
    .io_spriteVisible_9(gameLogic_io_spriteVisible_9),
    .io_spriteVisible_10(gameLogic_io_spriteVisible_10),
    .io_spriteVisible_11(gameLogic_io_spriteVisible_11),
    .io_spriteVisible_12(gameLogic_io_spriteVisible_12),
    .io_spriteVisible_13(gameLogic_io_spriteVisible_13),
    .io_spriteVisible_14(gameLogic_io_spriteVisible_14),
    .io_spriteVisible_15(gameLogic_io_spriteVisible_15),
    .io_spriteVisible_16(gameLogic_io_spriteVisible_16),
    .io_spriteVisible_17(gameLogic_io_spriteVisible_17),
    .io_spriteVisible_18(gameLogic_io_spriteVisible_18),
    .io_spriteVisible_19(gameLogic_io_spriteVisible_19),
    .io_spriteVisible_20(gameLogic_io_spriteVisible_20),
    .io_spriteVisible_21(gameLogic_io_spriteVisible_21),
    .io_spriteVisible_22(gameLogic_io_spriteVisible_22),
    .io_spriteVisible_23(gameLogic_io_spriteVisible_23),
    .io_spriteVisible_24(gameLogic_io_spriteVisible_24),
    .io_spriteVisible_25(gameLogic_io_spriteVisible_25),
    .io_spriteVisible_26(gameLogic_io_spriteVisible_26),
    .io_spriteVisible_27(gameLogic_io_spriteVisible_27),
    .io_spriteVisible_28(gameLogic_io_spriteVisible_28),
    .io_spriteVisible_29(gameLogic_io_spriteVisible_29),
    .io_spriteVisible_30(gameLogic_io_spriteVisible_30),
    .io_spriteVisible_31(gameLogic_io_spriteVisible_31),
    .io_spriteVisible_32(gameLogic_io_spriteVisible_32),
    .io_spriteVisible_33(gameLogic_io_spriteVisible_33),
    .io_spriteVisible_34(gameLogic_io_spriteVisible_34),
    .io_spriteVisible_35(gameLogic_io_spriteVisible_35),
    .io_spriteVisible_36(gameLogic_io_spriteVisible_36),
    .io_spriteVisible_37(gameLogic_io_spriteVisible_37),
    .io_spriteVisible_38(gameLogic_io_spriteVisible_38),
    .io_spriteVisible_39(gameLogic_io_spriteVisible_39),
    .io_spriteVisible_40(gameLogic_io_spriteVisible_40),
    .io_spriteVisible_41(gameLogic_io_spriteVisible_41),
    .io_spriteVisible_42(gameLogic_io_spriteVisible_42),
    .io_spriteVisible_43(gameLogic_io_spriteVisible_43),
    .io_spriteVisible_44(gameLogic_io_spriteVisible_44),
    .io_spriteVisible_45(gameLogic_io_spriteVisible_45),
    .io_spriteVisible_46(gameLogic_io_spriteVisible_46),
    .io_spriteVisible_47(gameLogic_io_spriteVisible_47),
    .io_spriteVisible_48(gameLogic_io_spriteVisible_48),
    .io_spriteVisible_49(gameLogic_io_spriteVisible_49),
    .io_spriteVisible_50(gameLogic_io_spriteVisible_50),
    .io_spriteVisible_51(gameLogic_io_spriteVisible_51),
    .io_spriteVisible_52(gameLogic_io_spriteVisible_52),
    .io_spriteVisible_53(gameLogic_io_spriteVisible_53),
    .io_spriteVisible_54(gameLogic_io_spriteVisible_54),
    .io_spriteVisible_55(gameLogic_io_spriteVisible_55),
    .io_spriteVisible_56(gameLogic_io_spriteVisible_56),
    .io_spriteVisible_57(gameLogic_io_spriteVisible_57),
    .io_spriteVisible_58(gameLogic_io_spriteVisible_58),
    .io_spriteVisible_59(gameLogic_io_spriteVisible_59),
    .io_spriteVisible_60(gameLogic_io_spriteVisible_60),
    .io_spriteVisible_61(gameLogic_io_spriteVisible_61),
    .io_spriteVisible_62(gameLogic_io_spriteVisible_62),
    .io_spriteVisible_63(gameLogic_io_spriteVisible_63),
    .io_spriteScaleUpHorizontal_16(gameLogic_io_spriteScaleUpHorizontal_16),
    .io_spriteScaleUpHorizontal_17(gameLogic_io_spriteScaleUpHorizontal_17),
    .io_spriteScaleUpHorizontal_18(gameLogic_io_spriteScaleUpHorizontal_18),
    .io_spriteScaleUpHorizontal_19(gameLogic_io_spriteScaleUpHorizontal_19),
    .io_spriteScaleUpHorizontal_20(gameLogic_io_spriteScaleUpHorizontal_20),
    .io_spriteScaleUpHorizontal_21(gameLogic_io_spriteScaleUpHorizontal_21),
    .io_spriteScaleUpHorizontal_22(gameLogic_io_spriteScaleUpHorizontal_22),
    .io_spriteScaleUpHorizontal_23(gameLogic_io_spriteScaleUpHorizontal_23),
    .io_spriteScaleUpHorizontal_24(gameLogic_io_spriteScaleUpHorizontal_24),
    .io_spriteScaleUpHorizontal_25(gameLogic_io_spriteScaleUpHorizontal_25),
    .io_spriteScaleUpHorizontal_26(gameLogic_io_spriteScaleUpHorizontal_26),
    .io_spriteScaleUpHorizontal_27(gameLogic_io_spriteScaleUpHorizontal_27),
    .io_spriteScaleUpHorizontal_28(gameLogic_io_spriteScaleUpHorizontal_28),
    .io_spriteScaleUpHorizontal_29(gameLogic_io_spriteScaleUpHorizontal_29),
    .io_spriteScaleUpHorizontal_30(gameLogic_io_spriteScaleUpHorizontal_30),
    .io_spriteScaleUpHorizontal_31(gameLogic_io_spriteScaleUpHorizontal_31),
    .io_spriteScaleUpHorizontal_32(gameLogic_io_spriteScaleUpHorizontal_32),
    .io_spriteScaleUpHorizontal_33(gameLogic_io_spriteScaleUpHorizontal_33),
    .io_spriteScaleUpHorizontal_34(gameLogic_io_spriteScaleUpHorizontal_34),
    .io_spriteScaleUpHorizontal_35(gameLogic_io_spriteScaleUpHorizontal_35),
    .io_spriteScaleUpHorizontal_36(gameLogic_io_spriteScaleUpHorizontal_36),
    .io_spriteScaleUpHorizontal_37(gameLogic_io_spriteScaleUpHorizontal_37),
    .io_spriteScaleUpHorizontal_38(gameLogic_io_spriteScaleUpHorizontal_38),
    .io_spriteScaleUpHorizontal_39(gameLogic_io_spriteScaleUpHorizontal_39),
    .io_spriteScaleUpHorizontal_40(gameLogic_io_spriteScaleUpHorizontal_40),
    .io_spriteScaleUpHorizontal_41(gameLogic_io_spriteScaleUpHorizontal_41),
    .io_spriteScaleUpHorizontal_42(gameLogic_io_spriteScaleUpHorizontal_42),
    .io_spriteScaleUpHorizontal_43(gameLogic_io_spriteScaleUpHorizontal_43),
    .io_spriteScaleUpHorizontal_44(gameLogic_io_spriteScaleUpHorizontal_44),
    .io_spriteScaleUpHorizontal_45(gameLogic_io_spriteScaleUpHorizontal_45),
    .io_spriteScaleUpHorizontal_58(gameLogic_io_spriteScaleUpHorizontal_58),
    .io_spriteScaleUpHorizontal_59(gameLogic_io_spriteScaleUpHorizontal_59),
    .io_spriteScaleUpHorizontal_60(gameLogic_io_spriteScaleUpHorizontal_60),
    .io_spriteScaleUpVertical_16(gameLogic_io_spriteScaleUpVertical_16),
    .io_spriteScaleUpVertical_17(gameLogic_io_spriteScaleUpVertical_17),
    .io_spriteScaleUpVertical_18(gameLogic_io_spriteScaleUpVertical_18),
    .io_spriteScaleUpVertical_19(gameLogic_io_spriteScaleUpVertical_19),
    .io_spriteScaleUpVertical_20(gameLogic_io_spriteScaleUpVertical_20),
    .io_spriteScaleUpVertical_21(gameLogic_io_spriteScaleUpVertical_21),
    .io_spriteScaleUpVertical_22(gameLogic_io_spriteScaleUpVertical_22),
    .io_spriteScaleUpVertical_23(gameLogic_io_spriteScaleUpVertical_23),
    .io_spriteScaleUpVertical_24(gameLogic_io_spriteScaleUpVertical_24),
    .io_spriteScaleUpVertical_25(gameLogic_io_spriteScaleUpVertical_25),
    .io_spriteScaleUpVertical_26(gameLogic_io_spriteScaleUpVertical_26),
    .io_spriteScaleUpVertical_27(gameLogic_io_spriteScaleUpVertical_27),
    .io_spriteScaleUpVertical_28(gameLogic_io_spriteScaleUpVertical_28),
    .io_spriteScaleUpVertical_29(gameLogic_io_spriteScaleUpVertical_29),
    .io_spriteScaleUpVertical_30(gameLogic_io_spriteScaleUpVertical_30),
    .io_spriteScaleUpVertical_31(gameLogic_io_spriteScaleUpVertical_31),
    .io_spriteScaleUpVertical_32(gameLogic_io_spriteScaleUpVertical_32),
    .io_spriteScaleUpVertical_33(gameLogic_io_spriteScaleUpVertical_33),
    .io_spriteScaleUpVertical_34(gameLogic_io_spriteScaleUpVertical_34),
    .io_spriteScaleUpVertical_35(gameLogic_io_spriteScaleUpVertical_35),
    .io_spriteScaleUpVertical_36(gameLogic_io_spriteScaleUpVertical_36),
    .io_spriteScaleUpVertical_37(gameLogic_io_spriteScaleUpVertical_37),
    .io_spriteScaleUpVertical_38(gameLogic_io_spriteScaleUpVertical_38),
    .io_spriteScaleUpVertical_39(gameLogic_io_spriteScaleUpVertical_39),
    .io_spriteScaleUpVertical_40(gameLogic_io_spriteScaleUpVertical_40),
    .io_spriteScaleUpVertical_41(gameLogic_io_spriteScaleUpVertical_41),
    .io_spriteScaleUpVertical_42(gameLogic_io_spriteScaleUpVertical_42),
    .io_spriteScaleUpVertical_43(gameLogic_io_spriteScaleUpVertical_43),
    .io_spriteScaleUpVertical_44(gameLogic_io_spriteScaleUpVertical_44),
    .io_spriteScaleUpVertical_45(gameLogic_io_spriteScaleUpVertical_45),
    .io_spriteScaleUpVertical_58(gameLogic_io_spriteScaleUpVertical_58),
    .io_spriteScaleUpVertical_59(gameLogic_io_spriteScaleUpVertical_59),
    .io_spriteScaleUpVertical_60(gameLogic_io_spriteScaleUpVertical_60),
    .io_viewBoxX(gameLogic_io_viewBoxX),
    .io_viewBoxY(gameLogic_io_viewBoxY),
    .io_newFrame(gameLogic_io_newFrame),
    .io_frameUpdateDone(gameLogic_io_frameUpdateDone)
  );
  assign io_vgaRed = graphicEngineVGA_io_vgaRed; // @[\\src\\main\\scala\\GameTop.scala 105:13]
  assign io_vgaBlue = graphicEngineVGA_io_vgaBlue; // @[\\src\\main\\scala\\GameTop.scala 107:14]
  assign io_vgaGreen = graphicEngineVGA_io_vgaGreen; // @[\\src\\main\\scala\\GameTop.scala 106:15]
  assign io_Hsync = graphicEngineVGA_io_Hsync; // @[\\src\\main\\scala\\GameTop.scala 108:12]
  assign io_Vsync = graphicEngineVGA_io_Vsync; // @[\\src\\main\\scala\\GameTop.scala 109:12]
  assign io_missingFrameError = graphicEngineVGA_io_missingFrameError; // @[\\src\\main\\scala\\GameTop.scala 120:24]
  assign io_viewBoxOutOfRangeError = graphicEngineVGA_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\GameTop.scala 122:29]
  assign graphicEngineVGA_clock = clock;
  assign graphicEngineVGA_reset = resetReleaseCounter == 22'h3d08ff ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameTop.scala 83:67 84:18 86:18]
  assign graphicEngineVGA_io_spriteXPosition_3 = gameLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_7 = gameLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_8 = gameLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_9 = gameLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_10 = gameLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_11 = gameLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_12 = gameLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_13 = gameLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_14 = gameLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_16 = gameLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_17 = gameLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_18 = gameLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_19 = gameLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_20 = gameLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_21 = gameLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_22 = gameLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_23 = gameLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_24 = gameLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_25 = gameLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_26 = gameLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_27 = gameLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_28 = gameLogic_io_spriteXPosition_28; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_29 = gameLogic_io_spriteXPosition_29; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_30 = gameLogic_io_spriteXPosition_30; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_31 = gameLogic_io_spriteXPosition_31; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_32 = gameLogic_io_spriteXPosition_32; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_33 = gameLogic_io_spriteXPosition_33; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_34 = gameLogic_io_spriteXPosition_34; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_35 = gameLogic_io_spriteXPosition_35; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_36 = gameLogic_io_spriteXPosition_36; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_37 = gameLogic_io_spriteXPosition_37; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_38 = gameLogic_io_spriteXPosition_38; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_39 = gameLogic_io_spriteXPosition_39; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_40 = gameLogic_io_spriteXPosition_40; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_41 = gameLogic_io_spriteXPosition_41; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_42 = gameLogic_io_spriteXPosition_42; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_43 = gameLogic_io_spriteXPosition_43; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_44 = gameLogic_io_spriteXPosition_44; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_45 = gameLogic_io_spriteXPosition_45; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_46 = gameLogic_io_spriteXPosition_46; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_47 = gameLogic_io_spriteXPosition_47; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_48 = gameLogic_io_spriteXPosition_48; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_49 = gameLogic_io_spriteXPosition_49; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_50 = gameLogic_io_spriteXPosition_50; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_51 = gameLogic_io_spriteXPosition_51; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_52 = gameLogic_io_spriteXPosition_52; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_53 = gameLogic_io_spriteXPosition_53; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_54 = gameLogic_io_spriteXPosition_54; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_55 = gameLogic_io_spriteXPosition_55; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_56 = gameLogic_io_spriteXPosition_56; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_57 = gameLogic_io_spriteXPosition_57; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_58 = gameLogic_io_spriteXPosition_58; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_59 = gameLogic_io_spriteXPosition_59; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_60 = gameLogic_io_spriteXPosition_60; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_61 = gameLogic_io_spriteXPosition_61; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_62 = gameLogic_io_spriteXPosition_62; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_63 = gameLogic_io_spriteXPosition_63; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteYPosition_3 = gameLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_7 = gameLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_8 = gameLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_9 = gameLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_10 = gameLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_11 = gameLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_12 = gameLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_13 = gameLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_14 = gameLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_16 = gameLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_17 = gameLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_18 = gameLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_19 = gameLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_20 = gameLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_21 = gameLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_22 = gameLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_23 = gameLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_24 = gameLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_25 = gameLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_26 = gameLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_27 = gameLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_28 = gameLogic_io_spriteYPosition_28; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_29 = gameLogic_io_spriteYPosition_29; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_30 = gameLogic_io_spriteYPosition_30; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_31 = gameLogic_io_spriteYPosition_31; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_32 = gameLogic_io_spriteYPosition_32; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_33 = gameLogic_io_spriteYPosition_33; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_34 = gameLogic_io_spriteYPosition_34; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_35 = gameLogic_io_spriteYPosition_35; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_36 = gameLogic_io_spriteYPosition_36; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_37 = gameLogic_io_spriteYPosition_37; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_38 = gameLogic_io_spriteYPosition_38; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_39 = gameLogic_io_spriteYPosition_39; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_40 = gameLogic_io_spriteYPosition_40; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_41 = gameLogic_io_spriteYPosition_41; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_42 = gameLogic_io_spriteYPosition_42; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_43 = gameLogic_io_spriteYPosition_43; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_44 = gameLogic_io_spriteYPosition_44; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_45 = gameLogic_io_spriteYPosition_45; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_46 = gameLogic_io_spriteYPosition_46; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_47 = gameLogic_io_spriteYPosition_47; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_48 = gameLogic_io_spriteYPosition_48; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_49 = gameLogic_io_spriteYPosition_49; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_50 = gameLogic_io_spriteYPosition_50; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_51 = gameLogic_io_spriteYPosition_51; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_52 = gameLogic_io_spriteYPosition_52; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_53 = gameLogic_io_spriteYPosition_53; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_54 = gameLogic_io_spriteYPosition_54; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_55 = gameLogic_io_spriteYPosition_55; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_56 = gameLogic_io_spriteYPosition_56; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_57 = gameLogic_io_spriteYPosition_57; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_58 = gameLogic_io_spriteYPosition_58; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_59 = gameLogic_io_spriteYPosition_59; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_60 = gameLogic_io_spriteYPosition_60; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_61 = gameLogic_io_spriteYPosition_61; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_62 = gameLogic_io_spriteYPosition_62; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_63 = gameLogic_io_spriteYPosition_63; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteVisible_3 = gameLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_4 = gameLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_5 = gameLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_6 = gameLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_7 = gameLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_8 = gameLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_9 = gameLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_10 = gameLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_11 = gameLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_12 = gameLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_13 = gameLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_14 = gameLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_15 = gameLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_16 = gameLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_17 = gameLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_18 = gameLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_19 = gameLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_20 = gameLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_21 = gameLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_22 = gameLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_23 = gameLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_24 = gameLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_25 = gameLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_26 = gameLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_27 = gameLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_28 = gameLogic_io_spriteVisible_28; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_29 = gameLogic_io_spriteVisible_29; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_30 = gameLogic_io_spriteVisible_30; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_31 = gameLogic_io_spriteVisible_31; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_32 = gameLogic_io_spriteVisible_32; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_33 = gameLogic_io_spriteVisible_33; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_34 = gameLogic_io_spriteVisible_34; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_35 = gameLogic_io_spriteVisible_35; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_36 = gameLogic_io_spriteVisible_36; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_37 = gameLogic_io_spriteVisible_37; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_38 = gameLogic_io_spriteVisible_38; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_39 = gameLogic_io_spriteVisible_39; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_40 = gameLogic_io_spriteVisible_40; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_41 = gameLogic_io_spriteVisible_41; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_42 = gameLogic_io_spriteVisible_42; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_43 = gameLogic_io_spriteVisible_43; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_44 = gameLogic_io_spriteVisible_44; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_45 = gameLogic_io_spriteVisible_45; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_46 = gameLogic_io_spriteVisible_46; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_47 = gameLogic_io_spriteVisible_47; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_48 = gameLogic_io_spriteVisible_48; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_49 = gameLogic_io_spriteVisible_49; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_50 = gameLogic_io_spriteVisible_50; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_51 = gameLogic_io_spriteVisible_51; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_52 = gameLogic_io_spriteVisible_52; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_53 = gameLogic_io_spriteVisible_53; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_54 = gameLogic_io_spriteVisible_54; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_55 = gameLogic_io_spriteVisible_55; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_56 = gameLogic_io_spriteVisible_56; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_57 = gameLogic_io_spriteVisible_57; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_58 = gameLogic_io_spriteVisible_58; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_59 = gameLogic_io_spriteVisible_59; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_60 = gameLogic_io_spriteVisible_60; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_61 = gameLogic_io_spriteVisible_61; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_62 = gameLogic_io_spriteVisible_62; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_63 = gameLogic_io_spriteVisible_63; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_16 = gameLogic_io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_17 = gameLogic_io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_18 = gameLogic_io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_19 = gameLogic_io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_20 = gameLogic_io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_21 = gameLogic_io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_22 = gameLogic_io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_23 = gameLogic_io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_24 = gameLogic_io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_25 = gameLogic_io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_26 = gameLogic_io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_27 = gameLogic_io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_28 = gameLogic_io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_29 = gameLogic_io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_30 = gameLogic_io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_31 = gameLogic_io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_32 = gameLogic_io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_33 = gameLogic_io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_34 = gameLogic_io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_35 = gameLogic_io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_36 = gameLogic_io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_37 = gameLogic_io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_38 = gameLogic_io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_39 = gameLogic_io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_40 = gameLogic_io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_41 = gameLogic_io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_42 = gameLogic_io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_43 = gameLogic_io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_44 = gameLogic_io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_45 = gameLogic_io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_58 = gameLogic_io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_59 = gameLogic_io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_60 = gameLogic_io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpVertical_16 = gameLogic_io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_17 = gameLogic_io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_18 = gameLogic_io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_19 = gameLogic_io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_20 = gameLogic_io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_21 = gameLogic_io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_22 = gameLogic_io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_23 = gameLogic_io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_24 = gameLogic_io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_25 = gameLogic_io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_26 = gameLogic_io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_27 = gameLogic_io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_28 = gameLogic_io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_29 = gameLogic_io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_30 = gameLogic_io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_31 = gameLogic_io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_32 = gameLogic_io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_33 = gameLogic_io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_34 = gameLogic_io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_35 = gameLogic_io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_36 = gameLogic_io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_37 = gameLogic_io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_38 = gameLogic_io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_39 = gameLogic_io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_40 = gameLogic_io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_41 = gameLogic_io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_42 = gameLogic_io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_43 = gameLogic_io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_44 = gameLogic_io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_45 = gameLogic_io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_58 = gameLogic_io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_59 = gameLogic_io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_60 = gameLogic_io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_viewBoxX = gameLogic_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 138:32]
  assign graphicEngineVGA_io_viewBoxY = gameLogic_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 139:32]
  assign graphicEngineVGA_io_frameUpdateDone = gameLogic_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 148:39]
  assign soundEngine_clock = clock;
  assign soundEngine_reset = reset;
  assign gameLogic_clock = clock;
  assign gameLogic_reset = resetReleaseCounter == 22'h3d08ff ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameTop.scala 83:67 84:18 86:18]
  assign gameLogic_io_btnC = btnCState; // @[\\src\\main\\scala\\GameTop.scala 98:21]
  assign gameLogic_io_btnU = btnUState; // @[\\src\\main\\scala\\GameTop.scala 99:21]
  assign gameLogic_io_btnL = btnLState; // @[\\src\\main\\scala\\GameTop.scala 100:21]
  assign gameLogic_io_btnR = btnRState; // @[\\src\\main\\scala\\GameTop.scala 101:21]
  assign gameLogic_io_btnD = btnDState; // @[\\src\\main\\scala\\GameTop.scala 102:21]
  assign gameLogic_io_newFrame = graphicEngineVGA_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 147:25]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 68:32]
      debounceCounter <= 21'h0; // @[\\src\\main\\scala\\GameTop.scala 68:32]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 70:57]
      debounceCounter <= 21'h0; // @[\\src\\main\\scala\\GameTop.scala 71:21]
    end else begin
      debounceCounter <= _debounceCounter_T_1; // @[\\src\\main\\scala\\GameTop.scala 74:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 81:36]
      resetReleaseCounter <= 22'h0; // @[\\src\\main\\scala\\GameTop.scala 81:36]
    end else if (!(resetReleaseCounter == 22'h3d08ff)) begin // @[\\src\\main\\scala\\GameTop.scala 83:67]
      resetReleaseCounter <= _resetReleaseCounter_T_1; // @[\\src\\main\\scala\\GameTop.scala 87:25]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnCState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnCState_pipeReg_0 <= btnCState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnCState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnCState_pipeReg_1 <= btnCState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnCState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnCState_pipeReg_2 <= io_btnC; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 93:28]
      btnCState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 93:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 93:28]
      btnCState <= btnCState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 93:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_0 <= btnUState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_1 <= btnUState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_2 <= io_btnU; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 94:28]
      btnUState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 94:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 94:28]
      btnUState <= btnUState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 94:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_0 <= btnLState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_1 <= btnLState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_2 <= io_btnL; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 95:28]
      btnLState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 95:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 95:28]
      btnLState <= btnLState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 95:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_0 <= btnRState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_1 <= btnRState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_2 <= io_btnR; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 96:28]
      btnRState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 96:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 96:28]
      btnRState <= btnRState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 96:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_0 <= btnDState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_1 <= btnDState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_2 <= io_btnD; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 97:28]
      btnDState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 97:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 97:28]
      btnDState <= btnDState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 97:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounceCounter = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  resetReleaseCounter = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btnCState_pipeReg_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  btnCState_pipeReg_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  btnCState_pipeReg_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  btnCState = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  btnUState_pipeReg_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  btnUState_pipeReg_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  btnUState_pipeReg_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btnUState = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  btnLState_pipeReg_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  btnLState_pipeReg_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  btnLState_pipeReg_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btnLState = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  btnRState_pipeReg_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  btnRState_pipeReg_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  btnRState_pipeReg_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  btnRState = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  btnDState_pipeReg_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  btnDState_pipeReg_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  btnDState_pipeReg_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  btnDState = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input        clock,
  input        reset,
  input        io_btnC, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnU, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnL, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnR, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnD, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaRed, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaGreen, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaBlue, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_Hsync, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_Vsync, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_0, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_1, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_2, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_3, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_4, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_5, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_6, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_7, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_0, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_1, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_2, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_3, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_4, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_5, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_6, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_7, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_missingFrameError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_backBufferWriteError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_viewBoxOutOfRangeError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_soundOut // @[\\src\\main\\scala\\Top.scala 14:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  gameTop_clock; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_reset; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnC; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnU; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnL; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnR; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnD; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaRed; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaBlue; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaGreen; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_Hsync; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_Vsync; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_missingFrameError; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\Top.scala 44:23]
  reg  syncResetInput_REG; // @[\\src\\main\\scala\\Top.scala 49:48]
  reg  syncResetInput_REG_1; // @[\\src\\main\\scala\\Top.scala 49:40]
  reg  syncResetInput_REG_2; // @[\\src\\main\\scala\\Top.scala 49:32]
  reg  pipeResetReg_0; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_1; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_2; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_3; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_4; // @[\\src\\main\\scala\\Top.scala 54:25]
  wire [4:0] _gameTop_reset_T = {pipeResetReg_4,pipeResetReg_3,pipeResetReg_2,pipeResetReg_1,pipeResetReg_0}; // @[\\src\\main\\scala\\Top.scala 59:33]
  GameTop gameTop ( // @[\\src\\main\\scala\\Top.scala 44:23]
    .clock(gameTop_clock),
    .reset(gameTop_reset),
    .io_btnC(gameTop_io_btnC),
    .io_btnU(gameTop_io_btnU),
    .io_btnL(gameTop_io_btnL),
    .io_btnR(gameTop_io_btnR),
    .io_btnD(gameTop_io_btnD),
    .io_vgaRed(gameTop_io_vgaRed),
    .io_vgaBlue(gameTop_io_vgaBlue),
    .io_vgaGreen(gameTop_io_vgaGreen),
    .io_Hsync(gameTop_io_Hsync),
    .io_Vsync(gameTop_io_Vsync),
    .io_missingFrameError(gameTop_io_missingFrameError),
    .io_viewBoxOutOfRangeError(gameTop_io_viewBoxOutOfRangeError)
  );
  assign io_vgaRed = gameTop_io_vgaRed; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_vgaGreen = gameTop_io_vgaGreen; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_vgaBlue = gameTop_io_vgaBlue; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_Hsync = gameTop_io_Hsync; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_Vsync = gameTop_io_Vsync; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_0 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_1 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_2 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_3 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_4 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_5 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_6 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_7 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_missingFrameError = gameTop_io_missingFrameError; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_backBufferWriteError = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_viewBoxOutOfRangeError = gameTop_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_soundOut = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_clock = clock;
  assign gameTop_reset = |_gameTop_reset_T; // @[\\src\\main\\scala\\Top.scala 59:40]
  assign gameTop_io_btnC = io_btnC; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnU = io_btnU; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnL = io_btnL; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnR = io_btnR; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnD = io_btnD; // @[\\src\\main\\scala\\Top.scala 62:14]
  always @(posedge clock) begin
    syncResetInput_REG <= reset; // @[\\src\\main\\scala\\Top.scala 49:48]
    syncResetInput_REG_1 <= syncResetInput_REG; // @[\\src\\main\\scala\\Top.scala 49:40]
    syncResetInput_REG_2 <= syncResetInput_REG_1; // @[\\src\\main\\scala\\Top.scala 49:32]
    pipeResetReg_0 <= pipeResetReg_1; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_1 <= pipeResetReg_2; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_2 <= pipeResetReg_3; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_3 <= pipeResetReg_4; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_4 <= ~syncResetInput_REG_2; // @[\\src\\main\\scala\\Top.scala 49:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  syncResetInput_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  syncResetInput_REG_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  syncResetInput_REG_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pipeResetReg_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pipeResetReg_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pipeResetReg_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pipeResetReg_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pipeResetReg_4 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
