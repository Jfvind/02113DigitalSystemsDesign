module Memory(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_1(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_2(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_2.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_3(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_3.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_4(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_4.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_5(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_5.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_6(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_6.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_7(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_7.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_8(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_8.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_9(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_9.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_10(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_10.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_11(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_11.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_12(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_12.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_13(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_13.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_14(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_14.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_15(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_15.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_16(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_16.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_17(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_17.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_18(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_18.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_19(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_19.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_20(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_20.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_21(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_21.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_22(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_22.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_23(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_23.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_24(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_24.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_25(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_25.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_26(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_26.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_27(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_27.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_28(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_28.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_29(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_29.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_30(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_30.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_31(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_31.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_32(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_32.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_33(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_33.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_34(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_34.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_35(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_35.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_36(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_36.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_37(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_37.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_38(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_38.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_39(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_39.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_40(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_40.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_41(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_41.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_42(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_42.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_43(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_43.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_44(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_44.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_45(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_45.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_46(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_46.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_47(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_47.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_48(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_48.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_49(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_49.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_50(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_50.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_51(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_51.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_52(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_52.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_53(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_53.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_54(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_54.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_55(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_55.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_56(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_56.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_57(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_57.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_58(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_58.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_59(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_59.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_60(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_60.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_61(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_61.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_62(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_62.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_63(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_63.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_64(
  input         clock,
  input  [10:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [5:0]  io_dataRead, // @[\\src\\main\\scala\\Memory.scala 48:14]
  input         io_writeEnable, // @[\\src\\main\\scala\\Memory.scala 48:14]
  input  [5:0]  io_dataWrite // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [10:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [5:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [5:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 57:26]
  RamSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(6)) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 57:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 63:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 58:21]
  assign ramsSpWf_we = io_writeEnable; // @[\\src\\main\\scala\\Memory.scala 59:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 60:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 61:22]
  assign ramsSpWf_di = io_dataWrite; // @[\\src\\main\\scala\\Memory.scala 62:20]
endmodule
module Memory_66(
  input         clock,
  input  [10:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [5:0]  io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [10:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [5:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [5:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(6), .LOAD_FILE("memory_init/backbuffer_init.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 6'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_67(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_68(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_69(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_2.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_70(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_3.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_71(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_4.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_72(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_5.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_73(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_6.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_74(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_7.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_75(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_8.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_76(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_9.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_77(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_10.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_78(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_11.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_79(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_12.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_80(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_13.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_81(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_14.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_82(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_15.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_83(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_16.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_84(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_17.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_85(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_18.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_86(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_19.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_87(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_20.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_88(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_21.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_89(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_22.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_90(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_23.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_91(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_24.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_92(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_25.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_93(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_26.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_94(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_27.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_95(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_28.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_96(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_29.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_97(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_30.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_98(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_31.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_99(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_32.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_100(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_33.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_101(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_34.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_102(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_35.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_103(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_36.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_104(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_37.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_105(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_38.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_106(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_39.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_107(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_40.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_108(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_41.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_109(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_42.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_110(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_43.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_111(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_44.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_112(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_45.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_113(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_46.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_114(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_47.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_115(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_48.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_116(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_49.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_117(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_50.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_118(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_51.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_119(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_52.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_120(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_53.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_121(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_54.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_122(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_55.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_123(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_56.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_124(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_57.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_125(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_58.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_126(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_59.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_127(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_60.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_128(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_61.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_129(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_62.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_130(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_63.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module MultiHotPriortyReductionTree(
  input  [5:0] io_dataInput_0, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_1, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_2, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_3, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_4, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_5, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_6, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_7, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_8, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_9, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_10, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_11, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_12, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_13, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_14, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_15, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_16, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_17, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_18, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_19, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_20, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_21, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_22, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_23, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_24, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_25, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_26, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_27, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_28, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_29, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_30, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_31, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_32, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_33, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_34, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_35, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_36, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_37, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_38, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_39, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_40, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_41, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_42, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_43, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_44, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_45, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_46, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_47, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_48, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_49, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_50, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_51, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_52, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_53, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_54, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_55, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_56, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_57, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_58, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_59, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_60, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_61, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_62, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_63, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_0, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_1, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_2, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_3, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_4, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_5, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_6, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_7, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_8, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_9, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_10, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_11, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_12, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_13, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_14, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_15, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_16, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_17, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_18, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_19, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_20, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_21, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_22, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_23, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_24, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_25, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_26, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_27, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_28, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_29, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_30, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_31, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_32, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_33, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_34, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_35, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_36, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_37, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_38, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_39, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_40, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_41, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_42, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_43, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_44, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_45, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_46, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_47, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_48, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_49, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_50, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_51, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_52, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_53, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_54, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_55, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_56, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_57, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_58, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_59, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_60, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_61, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_62, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_63, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  output [5:0] io_dataOutput, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  output       io_selectOutput // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
);
  wire  selectNodeOutputs_31 = io_selectInput_0 | io_selectInput_1; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_32 = io_selectInput_2 | io_selectInput_3; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_15 = selectNodeOutputs_31 | selectNodeOutputs_32; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_33 = io_selectInput_4 | io_selectInput_5; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_34 = io_selectInput_6 | io_selectInput_7; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_16 = selectNodeOutputs_33 | selectNodeOutputs_34; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_7 = selectNodeOutputs_15 | selectNodeOutputs_16; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_35 = io_selectInput_8 | io_selectInput_9; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_36 = io_selectInput_10 | io_selectInput_11; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_17 = selectNodeOutputs_35 | selectNodeOutputs_36; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_37 = io_selectInput_12 | io_selectInput_13; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_38 = io_selectInput_14 | io_selectInput_15; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_18 = selectNodeOutputs_37 | selectNodeOutputs_38; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_8 = selectNodeOutputs_17 | selectNodeOutputs_18; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_3 = selectNodeOutputs_7 | selectNodeOutputs_8; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_39 = io_selectInput_16 | io_selectInput_17; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_40 = io_selectInput_18 | io_selectInput_19; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_19 = selectNodeOutputs_39 | selectNodeOutputs_40; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_41 = io_selectInput_20 | io_selectInput_21; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_42 = io_selectInput_22 | io_selectInput_23; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_20 = selectNodeOutputs_41 | selectNodeOutputs_42; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_9 = selectNodeOutputs_19 | selectNodeOutputs_20; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_43 = io_selectInput_24 | io_selectInput_25; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_44 = io_selectInput_26 | io_selectInput_27; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_21 = selectNodeOutputs_43 | selectNodeOutputs_44; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_45 = io_selectInput_28 | io_selectInput_29; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_46 = io_selectInput_30 | io_selectInput_31; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_22 = selectNodeOutputs_45 | selectNodeOutputs_46; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_10 = selectNodeOutputs_21 | selectNodeOutputs_22; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_4 = selectNodeOutputs_9 | selectNodeOutputs_10; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_1 = selectNodeOutputs_3 | selectNodeOutputs_4; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_31 = io_selectInput_0 ? io_dataInput_0 : io_dataInput_1; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_32 = io_selectInput_2 ? io_dataInput_2 : io_dataInput_3; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_15 = selectNodeOutputs_31 ? dataNodeOutputs_31 : dataNodeOutputs_32; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_33 = io_selectInput_4 ? io_dataInput_4 : io_dataInput_5; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_34 = io_selectInput_6 ? io_dataInput_6 : io_dataInput_7; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_16 = selectNodeOutputs_33 ? dataNodeOutputs_33 : dataNodeOutputs_34; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_7 = selectNodeOutputs_15 ? dataNodeOutputs_15 : dataNodeOutputs_16; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_35 = io_selectInput_8 ? io_dataInput_8 : io_dataInput_9; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_36 = io_selectInput_10 ? io_dataInput_10 : io_dataInput_11; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_17 = selectNodeOutputs_35 ? dataNodeOutputs_35 : dataNodeOutputs_36; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_37 = io_selectInput_12 ? io_dataInput_12 : io_dataInput_13; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_38 = io_selectInput_14 ? io_dataInput_14 : io_dataInput_15; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_18 = selectNodeOutputs_37 ? dataNodeOutputs_37 : dataNodeOutputs_38; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_8 = selectNodeOutputs_17 ? dataNodeOutputs_17 : dataNodeOutputs_18; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_3 = selectNodeOutputs_7 ? dataNodeOutputs_7 : dataNodeOutputs_8; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_39 = io_selectInput_16 ? io_dataInput_16 : io_dataInput_17; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_40 = io_selectInput_18 ? io_dataInput_18 : io_dataInput_19; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_19 = selectNodeOutputs_39 ? dataNodeOutputs_39 : dataNodeOutputs_40; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_41 = io_selectInput_20 ? io_dataInput_20 : io_dataInput_21; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_42 = io_selectInput_22 ? io_dataInput_22 : io_dataInput_23; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_20 = selectNodeOutputs_41 ? dataNodeOutputs_41 : dataNodeOutputs_42; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_9 = selectNodeOutputs_19 ? dataNodeOutputs_19 : dataNodeOutputs_20; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_43 = io_selectInput_24 ? io_dataInput_24 : io_dataInput_25; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_44 = io_selectInput_26 ? io_dataInput_26 : io_dataInput_27; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_21 = selectNodeOutputs_43 ? dataNodeOutputs_43 : dataNodeOutputs_44; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_45 = io_selectInput_28 ? io_dataInput_28 : io_dataInput_29; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_46 = io_selectInput_30 ? io_dataInput_30 : io_dataInput_31; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_22 = selectNodeOutputs_45 ? dataNodeOutputs_45 : dataNodeOutputs_46; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_10 = selectNodeOutputs_21 ? dataNodeOutputs_21 : dataNodeOutputs_22; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_4 = selectNodeOutputs_9 ? dataNodeOutputs_9 : dataNodeOutputs_10; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_1 = selectNodeOutputs_3 ? dataNodeOutputs_3 : dataNodeOutputs_4; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_47 = io_selectInput_32 | io_selectInput_33; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_48 = io_selectInput_34 | io_selectInput_35; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_23 = selectNodeOutputs_47 | selectNodeOutputs_48; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_49 = io_selectInput_36 | io_selectInput_37; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_50 = io_selectInput_38 | io_selectInput_39; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_24 = selectNodeOutputs_49 | selectNodeOutputs_50; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_11 = selectNodeOutputs_23 | selectNodeOutputs_24; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_51 = io_selectInput_40 | io_selectInput_41; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_52 = io_selectInput_42 | io_selectInput_43; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_25 = selectNodeOutputs_51 | selectNodeOutputs_52; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_53 = io_selectInput_44 | io_selectInput_45; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_54 = io_selectInput_46 | io_selectInput_47; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_26 = selectNodeOutputs_53 | selectNodeOutputs_54; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_12 = selectNodeOutputs_25 | selectNodeOutputs_26; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_5 = selectNodeOutputs_11 | selectNodeOutputs_12; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_47 = io_selectInput_32 ? io_dataInput_32 : io_dataInput_33; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_48 = io_selectInput_34 ? io_dataInput_34 : io_dataInput_35; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_23 = selectNodeOutputs_47 ? dataNodeOutputs_47 : dataNodeOutputs_48; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_49 = io_selectInput_36 ? io_dataInput_36 : io_dataInput_37; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_50 = io_selectInput_38 ? io_dataInput_38 : io_dataInput_39; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_24 = selectNodeOutputs_49 ? dataNodeOutputs_49 : dataNodeOutputs_50; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_11 = selectNodeOutputs_23 ? dataNodeOutputs_23 : dataNodeOutputs_24; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_51 = io_selectInput_40 ? io_dataInput_40 : io_dataInput_41; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_52 = io_selectInput_42 ? io_dataInput_42 : io_dataInput_43; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_25 = selectNodeOutputs_51 ? dataNodeOutputs_51 : dataNodeOutputs_52; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_53 = io_selectInput_44 ? io_dataInput_44 : io_dataInput_45; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_54 = io_selectInput_46 ? io_dataInput_46 : io_dataInput_47; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_26 = selectNodeOutputs_53 ? dataNodeOutputs_53 : dataNodeOutputs_54; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_12 = selectNodeOutputs_25 ? dataNodeOutputs_25 : dataNodeOutputs_26; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_5 = selectNodeOutputs_11 ? dataNodeOutputs_11 : dataNodeOutputs_12; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_55 = io_selectInput_48 | io_selectInput_49; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_56 = io_selectInput_50 | io_selectInput_51; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_27 = selectNodeOutputs_55 | selectNodeOutputs_56; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_57 = io_selectInput_52 | io_selectInput_53; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_58 = io_selectInput_54 | io_selectInput_55; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_28 = selectNodeOutputs_57 | selectNodeOutputs_58; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_13 = selectNodeOutputs_27 | selectNodeOutputs_28; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_55 = io_selectInput_48 ? io_dataInput_48 : io_dataInput_49; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_56 = io_selectInput_50 ? io_dataInput_50 : io_dataInput_51; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_27 = selectNodeOutputs_55 ? dataNodeOutputs_55 : dataNodeOutputs_56; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_57 = io_selectInput_52 ? io_dataInput_52 : io_dataInput_53; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_58 = io_selectInput_54 ? io_dataInput_54 : io_dataInput_55; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_28 = selectNodeOutputs_57 ? dataNodeOutputs_57 : dataNodeOutputs_58; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_13 = selectNodeOutputs_27 ? dataNodeOutputs_27 : dataNodeOutputs_28; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_59 = io_selectInput_56 | io_selectInput_57; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_60 = io_selectInput_58 | io_selectInput_59; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_29 = selectNodeOutputs_59 | selectNodeOutputs_60; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_59 = io_selectInput_56 ? io_dataInput_56 : io_dataInput_57; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_60 = io_selectInput_58 ? io_dataInput_58 : io_dataInput_59; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_29 = selectNodeOutputs_59 ? dataNodeOutputs_59 : dataNodeOutputs_60; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_61 = io_selectInput_60 | io_selectInput_61; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_61 = io_selectInput_60 ? io_dataInput_60 : io_dataInput_61; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_62 = io_selectInput_62 ? io_dataInput_62 : io_dataInput_63; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_30 = selectNodeOutputs_61 ? dataNodeOutputs_61 : dataNodeOutputs_62; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_14 = selectNodeOutputs_29 ? dataNodeOutputs_29 : dataNodeOutputs_30; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_6 = selectNodeOutputs_13 ? dataNodeOutputs_13 : dataNodeOutputs_14; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_2 = selectNodeOutputs_5 ? dataNodeOutputs_5 : dataNodeOutputs_6; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_62 = io_selectInput_62 | io_selectInput_63; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_30 = selectNodeOutputs_61 | selectNodeOutputs_62; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_14 = selectNodeOutputs_29 | selectNodeOutputs_30; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_6 = selectNodeOutputs_13 | selectNodeOutputs_14; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_2 = selectNodeOutputs_5 | selectNodeOutputs_6; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  assign io_dataOutput = selectNodeOutputs_1 ? dataNodeOutputs_1 : dataNodeOutputs_2; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  assign io_selectOutput = selectNodeOutputs_1 | selectNodeOutputs_2; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
endmodule
module GraphicEngineVGA(
  input         clock,
  input         reset,
  input  [10:0] io_spriteXPosition_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_46, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_47, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_48, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_49, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_50, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_51, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_52, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_53, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_54, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_55, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_56, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_57, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_61, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_62, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_63, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_46, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_47, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_48, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_49, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_50, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_51, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_52, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_53, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_54, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_55, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_56, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_57, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_61, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_62, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_63, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_4, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_5, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_6, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_15, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_46, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_47, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_48, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_49, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_50, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_51, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_52, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_53, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_54, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_55, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_56, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_57, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_61, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_62, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_63, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpHorizontal_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_28, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_29, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_30, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_31, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_32, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_33, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_34, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_35, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_36, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_37, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_38, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_39, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_40, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_41, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_42, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_43, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_44, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_45, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_58, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_59, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteScaleUpVertical_60, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_viewBoxX, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [8:0]  io_viewBoxY, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_newFrame, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_frameUpdateDone, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_missingFrameError, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_viewBoxOutOfRangeError, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaRed, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaBlue, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaGreen, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_Hsync, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_Vsync // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
`endif // RANDOMIZE_REG_INIT
  wire  backTileMemories_0_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_0_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_1_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_1_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_2_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_2_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_3_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_3_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_4_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_4_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_5_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_5_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_6_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_6_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_7_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_7_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_8_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_8_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_9_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_9_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_10_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_10_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_11_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_11_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_12_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_12_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_13_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_13_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_14_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_14_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_15_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_15_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_16_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_16_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_17_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_17_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_18_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_18_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_19_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_19_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_20_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_20_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_21_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_21_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_22_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_22_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_23_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_23_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_24_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_24_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_25_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_25_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_26_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_26_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_27_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_27_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_28_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_28_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_29_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_29_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_30_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_30_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_31_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_31_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_32_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_32_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_32_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_33_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_33_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_33_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_34_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_34_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_34_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_35_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_35_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_35_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_36_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_36_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_36_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_37_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_37_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_37_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_38_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_38_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_38_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_39_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_39_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_39_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_40_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_40_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_40_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_41_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_41_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_41_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_42_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_42_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_42_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_43_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_43_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_43_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_44_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_44_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_44_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_45_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_45_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_45_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_46_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_46_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_46_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_47_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_47_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_47_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_48_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_48_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_48_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_49_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_49_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_49_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_50_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_50_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_50_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_51_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_51_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_51_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_52_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_52_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_52_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_53_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_53_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_53_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_54_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_54_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_54_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_55_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_55_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_55_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_56_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_56_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_56_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_57_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_57_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_57_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_58_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_58_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_58_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_59_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_59_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_59_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_60_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_60_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_60_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_61_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_61_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_61_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_62_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_62_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_62_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_63_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_63_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_63_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backBufferMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [10:0] backBufferMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [5:0] backBufferMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire  backBufferMemory_io_writeEnable; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [5:0] backBufferMemory_io_dataWrite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire  backBufferShadowMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [10:0] backBufferShadowMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [5:0] backBufferShadowMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire  backBufferShadowMemory_io_writeEnable; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [5:0] backBufferShadowMemory_io_dataWrite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire  backBufferRestoreMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire [10:0] backBufferRestoreMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire [5:0] backBufferRestoreMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire  spriteMemories_0_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_0_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_1_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_1_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_2_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_2_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_3_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_3_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_4_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_4_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_5_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_5_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_6_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_6_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_7_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_7_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_8_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_8_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_9_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_9_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_10_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_10_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_11_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_11_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_12_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_12_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_13_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_13_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_14_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_14_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_15_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_15_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_16_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_16_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_17_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_17_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_18_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_18_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_19_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_19_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_20_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_20_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_21_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_21_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_22_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_22_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_23_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_23_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_24_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_24_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_25_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_25_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_26_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_26_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_27_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_27_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_28_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_28_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_29_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_29_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_30_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_30_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_31_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_31_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_32_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_32_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_32_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_33_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_33_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_33_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_34_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_34_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_34_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_35_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_35_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_35_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_36_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_36_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_36_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_37_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_37_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_37_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_38_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_38_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_38_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_39_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_39_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_39_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_40_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_40_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_40_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_41_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_41_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_41_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_42_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_42_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_42_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_43_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_43_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_43_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_44_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_44_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_44_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_45_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_45_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_45_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_46_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_46_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_46_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_47_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_47_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_47_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_48_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_48_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_48_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_49_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_49_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_49_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_50_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_50_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_50_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_51_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_51_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_51_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_52_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_52_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_52_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_53_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_53_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_53_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_54_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_54_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_54_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_55_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_55_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_55_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_56_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_56_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_56_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_57_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_57_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_57_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_58_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_58_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_58_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_59_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_59_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_59_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_60_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_60_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_60_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_61_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_61_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_61_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_62_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_62_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_62_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_63_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_63_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_63_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  reg [1:0] ScaleCounterReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
  reg [9:0] CounterXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
  reg [9:0] CounterYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
  wire  _T_2 = CounterYReg == 10'h20c; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 78:26]
  wire [9:0] _CounterYReg_T_1 = CounterYReg + 10'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 82:38]
  wire [9:0] _GEN_0 = CounterYReg == 10'h20c ? 10'h0 : _CounterYReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 78:131 79:23 82:23]
  wire [9:0] _CounterXReg_T_1 = CounterXReg + 10'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 85:36]
  wire  _GEN_4 = CounterXReg == 10'h31f & _T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129 71:15]
  wire [1:0] _ScaleCounterReg_T_1 = ScaleCounterReg + 2'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 88:42]
  wire  _GEN_8 = ScaleCounterReg == 2'h3 & _GEN_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 71:15 74:52]
  reg [11:0] backMemoryRestoreCounter; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
  wire  restoreEnabled = backMemoryRestoreCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:33]
  wire  run = restoreEnabled ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:70 209:9 213:9]
  wire  Hsync = CounterXReg >= 10'h290 & CounterXReg < 10'h2f0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 92:79]
  wire  Vsync = CounterYReg >= 10'h1ea & CounterYReg < 10'h1ec; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 93:79]
  reg  io_Hsync_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg [20:0] frameClockCount; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
  wire [20:0] _frameClockCount_T_2 = frameClockCount + 21'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 105:92]
  wire  preDisplayArea = frameClockCount >= 21'h199a1b; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 106:40]
  reg [10:0] spriteXPositionReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [9:0] spriteYPositionReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg  spriteVisibleReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  wire  _GEN_141 = io_newFrame ? 1'h0 : spriteVisibleReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_142 = io_newFrame ? 1'h0 : spriteVisibleReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_143 = io_newFrame ? 1'h0 : spriteVisibleReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_144 = io_newFrame ? io_spriteVisible_3 : spriteVisibleReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_145 = io_newFrame ? io_spriteVisible_4 : spriteVisibleReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_146 = io_newFrame ? io_spriteVisible_5 : spriteVisibleReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_147 = io_newFrame ? io_spriteVisible_6 : spriteVisibleReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_148 = io_newFrame ? io_spriteVisible_7 : spriteVisibleReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_149 = io_newFrame ? io_spriteVisible_8 : spriteVisibleReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_150 = io_newFrame ? io_spriteVisible_9 : spriteVisibleReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_151 = io_newFrame ? io_spriteVisible_10 : spriteVisibleReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_152 = io_newFrame ? io_spriteVisible_11 : spriteVisibleReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_153 = io_newFrame ? io_spriteVisible_12 : spriteVisibleReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_154 = io_newFrame ? io_spriteVisible_13 : spriteVisibleReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_155 = io_newFrame ? io_spriteVisible_14 : spriteVisibleReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_156 = io_newFrame ? io_spriteVisible_15 : spriteVisibleReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_157 = io_newFrame ? io_spriteVisible_16 : spriteVisibleReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_158 = io_newFrame ? io_spriteVisible_17 : spriteVisibleReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_159 = io_newFrame ? io_spriteVisible_18 : spriteVisibleReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_160 = io_newFrame ? io_spriteVisible_19 : spriteVisibleReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_161 = io_newFrame ? io_spriteVisible_20 : spriteVisibleReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_162 = io_newFrame ? io_spriteVisible_21 : spriteVisibleReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_163 = io_newFrame ? io_spriteVisible_22 : spriteVisibleReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_164 = io_newFrame ? io_spriteVisible_23 : spriteVisibleReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_165 = io_newFrame ? io_spriteVisible_24 : spriteVisibleReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_166 = io_newFrame ? io_spriteVisible_25 : spriteVisibleReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_167 = io_newFrame ? io_spriteVisible_26 : spriteVisibleReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_168 = io_newFrame ? io_spriteVisible_27 : spriteVisibleReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_169 = io_newFrame ? io_spriteVisible_28 : spriteVisibleReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_170 = io_newFrame ? io_spriteVisible_29 : spriteVisibleReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_171 = io_newFrame ? io_spriteVisible_30 : spriteVisibleReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_172 = io_newFrame ? io_spriteVisible_31 : spriteVisibleReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_173 = io_newFrame ? io_spriteVisible_32 : spriteVisibleReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_174 = io_newFrame ? io_spriteVisible_33 : spriteVisibleReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_175 = io_newFrame ? io_spriteVisible_34 : spriteVisibleReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_176 = io_newFrame ? io_spriteVisible_35 : spriteVisibleReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_177 = io_newFrame ? io_spriteVisible_36 : spriteVisibleReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_178 = io_newFrame ? io_spriteVisible_37 : spriteVisibleReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_179 = io_newFrame ? io_spriteVisible_38 : spriteVisibleReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_180 = io_newFrame ? io_spriteVisible_39 : spriteVisibleReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_181 = io_newFrame ? io_spriteVisible_40 : spriteVisibleReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_182 = io_newFrame ? io_spriteVisible_41 : spriteVisibleReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_183 = io_newFrame ? io_spriteVisible_42 : spriteVisibleReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_184 = io_newFrame ? io_spriteVisible_43 : spriteVisibleReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_185 = io_newFrame ? io_spriteVisible_44 : spriteVisibleReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_186 = io_newFrame ? io_spriteVisible_45 : spriteVisibleReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_187 = io_newFrame ? io_spriteVisible_46 : spriteVisibleReg_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_188 = io_newFrame ? io_spriteVisible_47 : spriteVisibleReg_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_189 = io_newFrame ? io_spriteVisible_48 : spriteVisibleReg_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_190 = io_newFrame ? io_spriteVisible_49 : spriteVisibleReg_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_191 = io_newFrame ? io_spriteVisible_50 : spriteVisibleReg_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_192 = io_newFrame ? io_spriteVisible_51 : spriteVisibleReg_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_193 = io_newFrame ? io_spriteVisible_52 : spriteVisibleReg_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_194 = io_newFrame ? io_spriteVisible_53 : spriteVisibleReg_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_195 = io_newFrame ? io_spriteVisible_54 : spriteVisibleReg_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_196 = io_newFrame ? io_spriteVisible_55 : spriteVisibleReg_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_197 = io_newFrame ? io_spriteVisible_56 : spriteVisibleReg_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_198 = io_newFrame ? io_spriteVisible_57 : spriteVisibleReg_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_199 = io_newFrame ? io_spriteVisible_58 : spriteVisibleReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_200 = io_newFrame ? io_spriteVisible_59 : spriteVisibleReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_201 = io_newFrame ? io_spriteVisible_60 : spriteVisibleReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_202 = io_newFrame ? io_spriteVisible_61 : spriteVisibleReg_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_203 = io_newFrame ? io_spriteVisible_62 : spriteVisibleReg_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_204 = io_newFrame ? io_spriteVisible_63 : spriteVisibleReg_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  reg  spriteScaleUpHorizontalReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpHorizontalReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
  reg  spriteScaleUpVerticalReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg  spriteScaleUpVerticalReg_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
  reg [9:0] viewBoxXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
  reg [8:0] viewBoxYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
  reg  missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
  reg  viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
  wire [9:0] viewBoxXClipped = viewBoxXReg >= 10'h280 ? 10'h280 : viewBoxXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 137:28]
  wire [8:0] viewBoxYClipped = viewBoxYReg >= 9'h1e0 ? 9'h1e0 : viewBoxYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 138:28]
  wire [10:0] pixelXBack = CounterXReg + viewBoxXClipped; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 139:27]
  wire [9:0] _GEN_1692 = {{1'd0}, viewBoxYClipped}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 140:27]
  wire [10:0] pixelYBack = CounterYReg + _GEN_1692; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 140:27]
  wire  _GEN_591 = viewBoxXReg > 10'h280 | viewBoxYReg > 9'h1e0 | viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 141:51 142:31 130:42]
  reg  newFrameStikyReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
  wire  _GEN_592 = io_newFrame | newFrameStikyReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 148:21 149:22 147:33]
  reg  REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:16]
  wire  _GEN_594 = newFrameStikyReg & io_newFrame | missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 154:41 155:26 128:37]
  wire [10:0] _backTileMemories_0_io_address_T_2 = 6'h20 * pixelYBack[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:75]
  wire [10:0] _GEN_1693 = {{6'd0}, pixelXBack[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:62]
  wire [11:0] _backTileMemories_0_io_address_T_3 = _GEN_1693 + _backTileMemories_0_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:62]
  reg [6:0] backTileMemoryDataRead_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [11:0] backMemoryCopyCounter; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
  wire  _T_7 = backMemoryCopyCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 187:32]
  wire [11:0] _backMemoryCopyCounter_T_1 = backMemoryCopyCounter + 12'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 188:54]
  wire  copyEnabled = preDisplayArea & _T_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23 198:17]
  reg  copyEnabledReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 200:31]
  wire [11:0] _backMemoryRestoreCounter_T_1 = backMemoryRestoreCounter + 12'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 206:58]
  reg [10:0] backBufferShadowMemory_io_address_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:67]
  wire [10:0] _backBufferShadowMemory_io_address_T_2 = copyEnabled ? backMemoryCopyCounter[10:0] : 11'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:105]
  reg  backBufferShadowMemory_io_writeEnable_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:71]
  reg [10:0] backBufferMemory_io_address_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:61]
  wire [11:0] _backBufferMemory_io_address_T_3 = 6'h28 * pixelYBack[10:5]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:130]
  wire [11:0] _GEN_1757 = {{6'd0}, pixelXBack[10:5]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:117]
  wire [12:0] _backBufferMemory_io_address_T_4 = _GEN_1757 + _backBufferMemory_io_address_T_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:117]
  wire [12:0] _backBufferMemory_io_address_T_5 = copyEnabledReg ? {{2'd0}, backBufferMemory_io_address_REG} :
    _backBufferMemory_io_address_T_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:37]
  reg [5:0] fullBackgroundColor_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:56]
  wire [6:0] _GEN_605 = 6'h1 == fullBackgroundColor_REG ? backTileMemoryDataRead_1_REG : backTileMemoryDataRead_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_606 = 6'h2 == fullBackgroundColor_REG ? backTileMemoryDataRead_2_REG : _GEN_605; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_607 = 6'h3 == fullBackgroundColor_REG ? backTileMemoryDataRead_3_REG : _GEN_606; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_608 = 6'h4 == fullBackgroundColor_REG ? backTileMemoryDataRead_4_REG : _GEN_607; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_609 = 6'h5 == fullBackgroundColor_REG ? backTileMemoryDataRead_5_REG : _GEN_608; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_610 = 6'h6 == fullBackgroundColor_REG ? backTileMemoryDataRead_6_REG : _GEN_609; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_611 = 6'h7 == fullBackgroundColor_REG ? backTileMemoryDataRead_7_REG : _GEN_610; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_612 = 6'h8 == fullBackgroundColor_REG ? backTileMemoryDataRead_8_REG : _GEN_611; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_613 = 6'h9 == fullBackgroundColor_REG ? backTileMemoryDataRead_9_REG : _GEN_612; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_614 = 6'ha == fullBackgroundColor_REG ? backTileMemoryDataRead_10_REG : _GEN_613; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_615 = 6'hb == fullBackgroundColor_REG ? backTileMemoryDataRead_11_REG : _GEN_614; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_616 = 6'hc == fullBackgroundColor_REG ? backTileMemoryDataRead_12_REG : _GEN_615; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_617 = 6'hd == fullBackgroundColor_REG ? backTileMemoryDataRead_13_REG : _GEN_616; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_618 = 6'he == fullBackgroundColor_REG ? backTileMemoryDataRead_14_REG : _GEN_617; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_619 = 6'hf == fullBackgroundColor_REG ? backTileMemoryDataRead_15_REG : _GEN_618; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_620 = 6'h10 == fullBackgroundColor_REG ? backTileMemoryDataRead_16_REG : _GEN_619; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_621 = 6'h11 == fullBackgroundColor_REG ? backTileMemoryDataRead_17_REG : _GEN_620; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_622 = 6'h12 == fullBackgroundColor_REG ? backTileMemoryDataRead_18_REG : _GEN_621; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_623 = 6'h13 == fullBackgroundColor_REG ? backTileMemoryDataRead_19_REG : _GEN_622; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_624 = 6'h14 == fullBackgroundColor_REG ? backTileMemoryDataRead_20_REG : _GEN_623; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_625 = 6'h15 == fullBackgroundColor_REG ? backTileMemoryDataRead_21_REG : _GEN_624; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_626 = 6'h16 == fullBackgroundColor_REG ? backTileMemoryDataRead_22_REG : _GEN_625; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_627 = 6'h17 == fullBackgroundColor_REG ? backTileMemoryDataRead_23_REG : _GEN_626; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_628 = 6'h18 == fullBackgroundColor_REG ? backTileMemoryDataRead_24_REG : _GEN_627; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_629 = 6'h19 == fullBackgroundColor_REG ? backTileMemoryDataRead_25_REG : _GEN_628; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_630 = 6'h1a == fullBackgroundColor_REG ? backTileMemoryDataRead_26_REG : _GEN_629; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_631 = 6'h1b == fullBackgroundColor_REG ? backTileMemoryDataRead_27_REG : _GEN_630; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_632 = 6'h1c == fullBackgroundColor_REG ? backTileMemoryDataRead_28_REG : _GEN_631; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_633 = 6'h1d == fullBackgroundColor_REG ? backTileMemoryDataRead_29_REG : _GEN_632; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_634 = 6'h1e == fullBackgroundColor_REG ? backTileMemoryDataRead_30_REG : _GEN_633; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_635 = 6'h1f == fullBackgroundColor_REG ? backTileMemoryDataRead_31_REG : _GEN_634; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_636 = 6'h20 == fullBackgroundColor_REG ? backTileMemoryDataRead_32_REG : _GEN_635; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_637 = 6'h21 == fullBackgroundColor_REG ? backTileMemoryDataRead_33_REG : _GEN_636; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_638 = 6'h22 == fullBackgroundColor_REG ? backTileMemoryDataRead_34_REG : _GEN_637; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_639 = 6'h23 == fullBackgroundColor_REG ? backTileMemoryDataRead_35_REG : _GEN_638; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_640 = 6'h24 == fullBackgroundColor_REG ? backTileMemoryDataRead_36_REG : _GEN_639; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_641 = 6'h25 == fullBackgroundColor_REG ? backTileMemoryDataRead_37_REG : _GEN_640; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_642 = 6'h26 == fullBackgroundColor_REG ? backTileMemoryDataRead_38_REG : _GEN_641; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_643 = 6'h27 == fullBackgroundColor_REG ? backTileMemoryDataRead_39_REG : _GEN_642; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_644 = 6'h28 == fullBackgroundColor_REG ? backTileMemoryDataRead_40_REG : _GEN_643; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_645 = 6'h29 == fullBackgroundColor_REG ? backTileMemoryDataRead_41_REG : _GEN_644; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_646 = 6'h2a == fullBackgroundColor_REG ? backTileMemoryDataRead_42_REG : _GEN_645; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_647 = 6'h2b == fullBackgroundColor_REG ? backTileMemoryDataRead_43_REG : _GEN_646; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_648 = 6'h2c == fullBackgroundColor_REG ? backTileMemoryDataRead_44_REG : _GEN_647; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_649 = 6'h2d == fullBackgroundColor_REG ? backTileMemoryDataRead_45_REG : _GEN_648; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_650 = 6'h2e == fullBackgroundColor_REG ? backTileMemoryDataRead_46_REG : _GEN_649; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_651 = 6'h2f == fullBackgroundColor_REG ? backTileMemoryDataRead_47_REG : _GEN_650; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_652 = 6'h30 == fullBackgroundColor_REG ? backTileMemoryDataRead_48_REG : _GEN_651; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_653 = 6'h31 == fullBackgroundColor_REG ? backTileMemoryDataRead_49_REG : _GEN_652; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_654 = 6'h32 == fullBackgroundColor_REG ? backTileMemoryDataRead_50_REG : _GEN_653; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_655 = 6'h33 == fullBackgroundColor_REG ? backTileMemoryDataRead_51_REG : _GEN_654; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_656 = 6'h34 == fullBackgroundColor_REG ? backTileMemoryDataRead_52_REG : _GEN_655; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_657 = 6'h35 == fullBackgroundColor_REG ? backTileMemoryDataRead_53_REG : _GEN_656; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_658 = 6'h36 == fullBackgroundColor_REG ? backTileMemoryDataRead_54_REG : _GEN_657; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_659 = 6'h37 == fullBackgroundColor_REG ? backTileMemoryDataRead_55_REG : _GEN_658; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_660 = 6'h38 == fullBackgroundColor_REG ? backTileMemoryDataRead_56_REG : _GEN_659; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_661 = 6'h39 == fullBackgroundColor_REG ? backTileMemoryDataRead_57_REG : _GEN_660; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_662 = 6'h3a == fullBackgroundColor_REG ? backTileMemoryDataRead_58_REG : _GEN_661; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_663 = 6'h3b == fullBackgroundColor_REG ? backTileMemoryDataRead_59_REG : _GEN_662; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_664 = 6'h3c == fullBackgroundColor_REG ? backTileMemoryDataRead_60_REG : _GEN_663; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_665 = 6'h3d == fullBackgroundColor_REG ? backTileMemoryDataRead_61_REG : _GEN_664; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_666 = 6'h3e == fullBackgroundColor_REG ? backTileMemoryDataRead_62_REG : _GEN_665; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] fullBackgroundColor = 6'h3f == fullBackgroundColor_REG ? backTileMemoryDataRead_63_REG : _GEN_666; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  reg [5:0] pixelColorBack; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 245:31]
  wire [10:0] _inSpriteXValue_T_1 = {1'h0,CounterXReg}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:47]
  wire [11:0] inSpriteXValue = $signed(_inSpriteXValue_T_1) - 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_0 = $signed(inSpriteXValue) >= 12'sh0 & $signed(inSpriteXValue) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_674 = {{1{inSpriteXValue[11]}},inSpriteXValue}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _inSpriteYValue_T_1 = {1'h0,CounterYReg}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:47]
  wire [11:0] inSpriteYValue = $signed(_inSpriteYValue_T_1) - 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_0 = inSpriteYValue[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_0 = $signed(inSpriteYPreScaled_0) >= 11'sh0 & $signed(inSpriteYPreScaled_0) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_682 = {{1{inSpriteYPreScaled_0[10]}},inSpriteYPreScaled_0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_3 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_3); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_3 = $signed(inSpriteXValue_3) >= 12'sh0 & $signed(inSpriteXValue_3) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_722 = {{1{inSpriteXValue_3[11]}},inSpriteXValue_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1761 = {{1{spriteYPositionReg_3[9]}},spriteYPositionReg_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_3 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1761); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_3 = inSpriteYValue_3[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_3 = $signed(inSpriteYPreScaled_3) >= 11'sh0 & $signed(inSpriteYPreScaled_3) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_730 = {{1{inSpriteYPreScaled_3[10]}},inSpriteYPreScaled_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_7 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_7); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_7 = $signed(inSpriteXValue_7) >= 12'sh0 & $signed(inSpriteXValue_7) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_786 = {{1{inSpriteXValue_7[11]}},inSpriteXValue_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1766 = {{1{spriteYPositionReg_7[9]}},spriteYPositionReg_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_7 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1766); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_7 = inSpriteYValue_7[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_7 = $signed(inSpriteYPreScaled_7) >= 11'sh0 & $signed(inSpriteYPreScaled_7) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_794 = {{1{inSpriteYPreScaled_7[10]}},inSpriteYPreScaled_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_8 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_8); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_8 = $signed(inSpriteXValue_8) >= 12'sh0 & $signed(inSpriteXValue_8) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_802 = {{1{inSpriteXValue_8[11]}},inSpriteXValue_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1768 = {{1{spriteYPositionReg_8[9]}},spriteYPositionReg_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_8 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1768); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_8 = inSpriteYValue_8[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_8 = $signed(inSpriteYPreScaled_8) >= 11'sh0 & $signed(inSpriteYPreScaled_8) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_810 = {{1{inSpriteYPreScaled_8[10]}},inSpriteYPreScaled_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_9 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_9); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_9 = $signed(inSpriteXValue_9) >= 12'sh0 & $signed(inSpriteXValue_9) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_818 = {{1{inSpriteXValue_9[11]}},inSpriteXValue_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1770 = {{1{spriteYPositionReg_9[9]}},spriteYPositionReg_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_9 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1770); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_9 = inSpriteYValue_9[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_9 = $signed(inSpriteYPreScaled_9) >= 11'sh0 & $signed(inSpriteYPreScaled_9) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_826 = {{1{inSpriteYPreScaled_9[10]}},inSpriteYPreScaled_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_10 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_10); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_10 = $signed(inSpriteXValue_10) >= 12'sh0 & $signed(inSpriteXValue_10) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_834 = {{1{inSpriteXValue_10[11]}},inSpriteXValue_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1772 = {{1{spriteYPositionReg_10[9]}},spriteYPositionReg_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_10 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1772); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_10 = inSpriteYValue_10[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_10 = $signed(inSpriteYPreScaled_10) >= 11'sh0 & $signed(inSpriteYPreScaled_10) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_842 = {{1{inSpriteYPreScaled_10[10]}},inSpriteYPreScaled_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_11 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_11); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_11 = $signed(inSpriteXValue_11) >= 12'sh0 & $signed(inSpriteXValue_11) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_850 = {{1{inSpriteXValue_11[11]}},inSpriteXValue_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1774 = {{1{spriteYPositionReg_11[9]}},spriteYPositionReg_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_11 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1774); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_11 = inSpriteYValue_11[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_11 = $signed(inSpriteYPreScaled_11) >= 11'sh0 & $signed(inSpriteYPreScaled_11) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_858 = {{1{inSpriteYPreScaled_11[10]}},inSpriteYPreScaled_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_12 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_12); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_12 = $signed(inSpriteXValue_12) >= 12'sh0 & $signed(inSpriteXValue_12) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_866 = {{1{inSpriteXValue_12[11]}},inSpriteXValue_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1776 = {{1{spriteYPositionReg_12[9]}},spriteYPositionReg_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_12 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1776); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_12 = inSpriteYValue_12[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_12 = $signed(inSpriteYPreScaled_12) >= 11'sh0 & $signed(inSpriteYPreScaled_12) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_874 = {{1{inSpriteYPreScaled_12[10]}},inSpriteYPreScaled_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_13 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_13); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_13 = $signed(inSpriteXValue_13) >= 12'sh0 & $signed(inSpriteXValue_13) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_882 = {{1{inSpriteXValue_13[11]}},inSpriteXValue_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1778 = {{1{spriteYPositionReg_13[9]}},spriteYPositionReg_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_13 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1778); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_13 = inSpriteYValue_13[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_13 = $signed(inSpriteYPreScaled_13) >= 11'sh0 & $signed(inSpriteYPreScaled_13) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_890 = {{1{inSpriteYPreScaled_13[10]}},inSpriteYPreScaled_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_14 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_14); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_14 = $signed(inSpriteXValue_14) >= 12'sh0 & $signed(inSpriteXValue_14) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_898 = {{1{inSpriteXValue_14[11]}},inSpriteXValue_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1780 = {{1{spriteYPositionReg_14[9]}},spriteYPositionReg_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_14 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1780); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_14 = inSpriteYValue_14[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_14 = $signed(inSpriteYPreScaled_14) >= 11'sh0 & $signed(inSpriteYPreScaled_14) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_906 = {{1{inSpriteYPreScaled_14[10]}},inSpriteYPreScaled_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_16 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_16); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_16_T = $signed(inSpriteXValue_16) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_16_T_4 = inSpriteXValue_16[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_16_T_8 = _inSpriteHorizontal_16_T & $signed(inSpriteXValue_16) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_16_T_5 = {$signed(inSpriteXValue_16), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_16_T_14 = _inSpriteHorizontal_16_T & $signed(inSpriteXValue_16) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_928 = spriteScaleUpHorizontalReg_16 ? $signed({{2{_inSpriteX_16_T_4[10]}},_inSpriteX_16_T_4}) :
    $signed(_inSpriteX_16_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_929 = spriteScaleUpHorizontalReg_16 ? _inSpriteHorizontal_16_T_8 : _inSpriteHorizontal_16_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_930 = ~spriteScaleUpHorizontalReg_16 ? $signed({{1{inSpriteXValue_16[11]}},inSpriteXValue_16}) :
    $signed(_GEN_928); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_16 = ~spriteScaleUpHorizontalReg_16 ? $signed(inSpriteXValue_16) >= 12'sh0 & $signed(
    inSpriteXValue_16) < 12'sh20 : _GEN_929; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1783 = {{1{spriteYPositionReg_16[9]}},spriteYPositionReg_16}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_16 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1783); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_16 = inSpriteYValue_16[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_16_T = $signed(inSpriteYPreScaled_16) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_16_T_4 = inSpriteYPreScaled_16[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_16_T_8 = _inSpriteVertical_16_T & $signed(inSpriteYPreScaled_16) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_16_T_5 = {$signed(inSpriteYPreScaled_16), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_16_T_14 = _inSpriteVertical_16_T & $signed(inSpriteYPreScaled_16) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_936 = spriteScaleUpVerticalReg_16 ? $signed({{2{_inSpriteY_16_T_4[9]}},_inSpriteY_16_T_4}) : $signed(
    _inSpriteY_16_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_937 = spriteScaleUpVerticalReg_16 ? _inSpriteVertical_16_T_8 : _inSpriteVertical_16_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_938 = ~spriteScaleUpVerticalReg_16 ? $signed({{1{inSpriteYPreScaled_16[10]}},inSpriteYPreScaled_16})
     : $signed(_GEN_936); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_16 = ~spriteScaleUpVerticalReg_16 ? $signed(inSpriteYPreScaled_16) >= 11'sh0 & $signed(
    inSpriteYPreScaled_16) < 11'sh20 : _GEN_937; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_17 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_17); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_17_T = $signed(inSpriteXValue_17) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_17_T_4 = inSpriteXValue_17[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_17_T_8 = _inSpriteHorizontal_17_T & $signed(inSpriteXValue_17) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_17_T_5 = {$signed(inSpriteXValue_17), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_17_T_14 = _inSpriteHorizontal_17_T & $signed(inSpriteXValue_17) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_944 = spriteScaleUpHorizontalReg_17 ? $signed({{2{_inSpriteX_17_T_4[10]}},_inSpriteX_17_T_4}) :
    $signed(_inSpriteX_17_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_945 = spriteScaleUpHorizontalReg_17 ? _inSpriteHorizontal_17_T_8 : _inSpriteHorizontal_17_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_946 = ~spriteScaleUpHorizontalReg_17 ? $signed({{1{inSpriteXValue_17[11]}},inSpriteXValue_17}) :
    $signed(_GEN_944); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_17 = ~spriteScaleUpHorizontalReg_17 ? $signed(inSpriteXValue_17) >= 12'sh0 & $signed(
    inSpriteXValue_17) < 12'sh20 : _GEN_945; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1785 = {{1{spriteYPositionReg_17[9]}},spriteYPositionReg_17}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_17 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1785); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_17 = inSpriteYValue_17[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_17_T = $signed(inSpriteYPreScaled_17) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_17_T_4 = inSpriteYPreScaled_17[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_17_T_8 = _inSpriteVertical_17_T & $signed(inSpriteYPreScaled_17) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_17_T_5 = {$signed(inSpriteYPreScaled_17), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_17_T_14 = _inSpriteVertical_17_T & $signed(inSpriteYPreScaled_17) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_952 = spriteScaleUpVerticalReg_17 ? $signed({{2{_inSpriteY_17_T_4[9]}},_inSpriteY_17_T_4}) : $signed(
    _inSpriteY_17_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_953 = spriteScaleUpVerticalReg_17 ? _inSpriteVertical_17_T_8 : _inSpriteVertical_17_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_954 = ~spriteScaleUpVerticalReg_17 ? $signed({{1{inSpriteYPreScaled_17[10]}},inSpriteYPreScaled_17})
     : $signed(_GEN_952); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_17 = ~spriteScaleUpVerticalReg_17 ? $signed(inSpriteYPreScaled_17) >= 11'sh0 & $signed(
    inSpriteYPreScaled_17) < 11'sh20 : _GEN_953; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_18 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_18); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_18_T = $signed(inSpriteXValue_18) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_18_T_4 = inSpriteXValue_18[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_18_T_8 = _inSpriteHorizontal_18_T & $signed(inSpriteXValue_18) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_18_T_5 = {$signed(inSpriteXValue_18), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_18_T_14 = _inSpriteHorizontal_18_T & $signed(inSpriteXValue_18) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_960 = spriteScaleUpHorizontalReg_18 ? $signed({{2{_inSpriteX_18_T_4[10]}},_inSpriteX_18_T_4}) :
    $signed(_inSpriteX_18_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_961 = spriteScaleUpHorizontalReg_18 ? _inSpriteHorizontal_18_T_8 : _inSpriteHorizontal_18_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_962 = ~spriteScaleUpHorizontalReg_18 ? $signed({{1{inSpriteXValue_18[11]}},inSpriteXValue_18}) :
    $signed(_GEN_960); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_18 = ~spriteScaleUpHorizontalReg_18 ? $signed(inSpriteXValue_18) >= 12'sh0 & $signed(
    inSpriteXValue_18) < 12'sh20 : _GEN_961; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1787 = {{1{spriteYPositionReg_18[9]}},spriteYPositionReg_18}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_18 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1787); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_18 = inSpriteYValue_18[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_18_T = $signed(inSpriteYPreScaled_18) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_18_T_4 = inSpriteYPreScaled_18[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_18_T_8 = _inSpriteVertical_18_T & $signed(inSpriteYPreScaled_18) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_18_T_5 = {$signed(inSpriteYPreScaled_18), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_18_T_14 = _inSpriteVertical_18_T & $signed(inSpriteYPreScaled_18) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_968 = spriteScaleUpVerticalReg_18 ? $signed({{2{_inSpriteY_18_T_4[9]}},_inSpriteY_18_T_4}) : $signed(
    _inSpriteY_18_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_969 = spriteScaleUpVerticalReg_18 ? _inSpriteVertical_18_T_8 : _inSpriteVertical_18_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_970 = ~spriteScaleUpVerticalReg_18 ? $signed({{1{inSpriteYPreScaled_18[10]}},inSpriteYPreScaled_18})
     : $signed(_GEN_968); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_18 = ~spriteScaleUpVerticalReg_18 ? $signed(inSpriteYPreScaled_18) >= 11'sh0 & $signed(
    inSpriteYPreScaled_18) < 11'sh20 : _GEN_969; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_19 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_19); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_19_T = $signed(inSpriteXValue_19) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_19_T_4 = inSpriteXValue_19[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_19_T_8 = _inSpriteHorizontal_19_T & $signed(inSpriteXValue_19) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_19_T_5 = {$signed(inSpriteXValue_19), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_19_T_14 = _inSpriteHorizontal_19_T & $signed(inSpriteXValue_19) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_976 = spriteScaleUpHorizontalReg_19 ? $signed({{2{_inSpriteX_19_T_4[10]}},_inSpriteX_19_T_4}) :
    $signed(_inSpriteX_19_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_977 = spriteScaleUpHorizontalReg_19 ? _inSpriteHorizontal_19_T_8 : _inSpriteHorizontal_19_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_978 = ~spriteScaleUpHorizontalReg_19 ? $signed({{1{inSpriteXValue_19[11]}},inSpriteXValue_19}) :
    $signed(_GEN_976); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_19 = ~spriteScaleUpHorizontalReg_19 ? $signed(inSpriteXValue_19) >= 12'sh0 & $signed(
    inSpriteXValue_19) < 12'sh20 : _GEN_977; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1789 = {{1{spriteYPositionReg_19[9]}},spriteYPositionReg_19}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_19 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1789); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_19 = inSpriteYValue_19[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_19_T = $signed(inSpriteYPreScaled_19) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_19_T_4 = inSpriteYPreScaled_19[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_19_T_8 = _inSpriteVertical_19_T & $signed(inSpriteYPreScaled_19) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_19_T_5 = {$signed(inSpriteYPreScaled_19), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_19_T_14 = _inSpriteVertical_19_T & $signed(inSpriteYPreScaled_19) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_984 = spriteScaleUpVerticalReg_19 ? $signed({{2{_inSpriteY_19_T_4[9]}},_inSpriteY_19_T_4}) : $signed(
    _inSpriteY_19_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_985 = spriteScaleUpVerticalReg_19 ? _inSpriteVertical_19_T_8 : _inSpriteVertical_19_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_986 = ~spriteScaleUpVerticalReg_19 ? $signed({{1{inSpriteYPreScaled_19[10]}},inSpriteYPreScaled_19})
     : $signed(_GEN_984); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_19 = ~spriteScaleUpVerticalReg_19 ? $signed(inSpriteYPreScaled_19) >= 11'sh0 & $signed(
    inSpriteYPreScaled_19) < 11'sh20 : _GEN_985; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_20 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_20); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_20_T = $signed(inSpriteXValue_20) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_20_T_4 = inSpriteXValue_20[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_20_T_8 = _inSpriteHorizontal_20_T & $signed(inSpriteXValue_20) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_20_T_5 = {$signed(inSpriteXValue_20), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_20_T_14 = _inSpriteHorizontal_20_T & $signed(inSpriteXValue_20) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_992 = spriteScaleUpHorizontalReg_20 ? $signed({{2{_inSpriteX_20_T_4[10]}},_inSpriteX_20_T_4}) :
    $signed(_inSpriteX_20_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_993 = spriteScaleUpHorizontalReg_20 ? _inSpriteHorizontal_20_T_8 : _inSpriteHorizontal_20_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_994 = ~spriteScaleUpHorizontalReg_20 ? $signed({{1{inSpriteXValue_20[11]}},inSpriteXValue_20}) :
    $signed(_GEN_992); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_20 = ~spriteScaleUpHorizontalReg_20 ? $signed(inSpriteXValue_20) >= 12'sh0 & $signed(
    inSpriteXValue_20) < 12'sh20 : _GEN_993; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1791 = {{1{spriteYPositionReg_20[9]}},spriteYPositionReg_20}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_20 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1791); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_20 = inSpriteYValue_20[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_20_T = $signed(inSpriteYPreScaled_20) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_20_T_4 = inSpriteYPreScaled_20[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_20_T_8 = _inSpriteVertical_20_T & $signed(inSpriteYPreScaled_20) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_20_T_5 = {$signed(inSpriteYPreScaled_20), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_20_T_14 = _inSpriteVertical_20_T & $signed(inSpriteYPreScaled_20) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1000 = spriteScaleUpVerticalReg_20 ? $signed({{2{_inSpriteY_20_T_4[9]}},_inSpriteY_20_T_4}) :
    $signed(_inSpriteY_20_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1001 = spriteScaleUpVerticalReg_20 ? _inSpriteVertical_20_T_8 : _inSpriteVertical_20_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1002 = ~spriteScaleUpVerticalReg_20 ? $signed({{1{inSpriteYPreScaled_20[10]}},inSpriteYPreScaled_20})
     : $signed(_GEN_1000); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_20 = ~spriteScaleUpVerticalReg_20 ? $signed(inSpriteYPreScaled_20) >= 11'sh0 & $signed(
    inSpriteYPreScaled_20) < 11'sh20 : _GEN_1001; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_21 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_21); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_21_T = $signed(inSpriteXValue_21) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_21_T_4 = inSpriteXValue_21[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_21_T_8 = _inSpriteHorizontal_21_T & $signed(inSpriteXValue_21) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_21_T_5 = {$signed(inSpriteXValue_21), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_21_T_14 = _inSpriteHorizontal_21_T & $signed(inSpriteXValue_21) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1008 = spriteScaleUpHorizontalReg_21 ? $signed({{2{_inSpriteX_21_T_4[10]}},_inSpriteX_21_T_4}) :
    $signed(_inSpriteX_21_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1009 = spriteScaleUpHorizontalReg_21 ? _inSpriteHorizontal_21_T_8 : _inSpriteHorizontal_21_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1010 = ~spriteScaleUpHorizontalReg_21 ? $signed({{1{inSpriteXValue_21[11]}},inSpriteXValue_21}) :
    $signed(_GEN_1008); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_21 = ~spriteScaleUpHorizontalReg_21 ? $signed(inSpriteXValue_21) >= 12'sh0 & $signed(
    inSpriteXValue_21) < 12'sh20 : _GEN_1009; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1793 = {{1{spriteYPositionReg_21[9]}},spriteYPositionReg_21}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_21 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1793); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_21 = inSpriteYValue_21[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_21_T = $signed(inSpriteYPreScaled_21) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_21_T_4 = inSpriteYPreScaled_21[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_21_T_8 = _inSpriteVertical_21_T & $signed(inSpriteYPreScaled_21) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_21_T_5 = {$signed(inSpriteYPreScaled_21), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_21_T_14 = _inSpriteVertical_21_T & $signed(inSpriteYPreScaled_21) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1016 = spriteScaleUpVerticalReg_21 ? $signed({{2{_inSpriteY_21_T_4[9]}},_inSpriteY_21_T_4}) :
    $signed(_inSpriteY_21_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1017 = spriteScaleUpVerticalReg_21 ? _inSpriteVertical_21_T_8 : _inSpriteVertical_21_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1018 = ~spriteScaleUpVerticalReg_21 ? $signed({{1{inSpriteYPreScaled_21[10]}},inSpriteYPreScaled_21})
     : $signed(_GEN_1016); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_21 = ~spriteScaleUpVerticalReg_21 ? $signed(inSpriteYPreScaled_21) >= 11'sh0 & $signed(
    inSpriteYPreScaled_21) < 11'sh20 : _GEN_1017; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_22 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_22); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_22_T = $signed(inSpriteXValue_22) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_22_T_4 = inSpriteXValue_22[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_22_T_8 = _inSpriteHorizontal_22_T & $signed(inSpriteXValue_22) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_22_T_5 = {$signed(inSpriteXValue_22), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_22_T_14 = _inSpriteHorizontal_22_T & $signed(inSpriteXValue_22) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1024 = spriteScaleUpHorizontalReg_22 ? $signed({{2{_inSpriteX_22_T_4[10]}},_inSpriteX_22_T_4}) :
    $signed(_inSpriteX_22_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1025 = spriteScaleUpHorizontalReg_22 ? _inSpriteHorizontal_22_T_8 : _inSpriteHorizontal_22_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1026 = ~spriteScaleUpHorizontalReg_22 ? $signed({{1{inSpriteXValue_22[11]}},inSpriteXValue_22}) :
    $signed(_GEN_1024); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_22 = ~spriteScaleUpHorizontalReg_22 ? $signed(inSpriteXValue_22) >= 12'sh0 & $signed(
    inSpriteXValue_22) < 12'sh20 : _GEN_1025; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1795 = {{1{spriteYPositionReg_22[9]}},spriteYPositionReg_22}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_22 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1795); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_22 = inSpriteYValue_22[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_22_T = $signed(inSpriteYPreScaled_22) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_22_T_4 = inSpriteYPreScaled_22[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_22_T_8 = _inSpriteVertical_22_T & $signed(inSpriteYPreScaled_22) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_22_T_5 = {$signed(inSpriteYPreScaled_22), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_22_T_14 = _inSpriteVertical_22_T & $signed(inSpriteYPreScaled_22) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1032 = spriteScaleUpVerticalReg_22 ? $signed({{2{_inSpriteY_22_T_4[9]}},_inSpriteY_22_T_4}) :
    $signed(_inSpriteY_22_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1033 = spriteScaleUpVerticalReg_22 ? _inSpriteVertical_22_T_8 : _inSpriteVertical_22_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1034 = ~spriteScaleUpVerticalReg_22 ? $signed({{1{inSpriteYPreScaled_22[10]}},inSpriteYPreScaled_22})
     : $signed(_GEN_1032); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_22 = ~spriteScaleUpVerticalReg_22 ? $signed(inSpriteYPreScaled_22) >= 11'sh0 & $signed(
    inSpriteYPreScaled_22) < 11'sh20 : _GEN_1033; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_23 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_23); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_23_T = $signed(inSpriteXValue_23) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_23_T_4 = inSpriteXValue_23[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_23_T_8 = _inSpriteHorizontal_23_T & $signed(inSpriteXValue_23) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_23_T_5 = {$signed(inSpriteXValue_23), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_23_T_14 = _inSpriteHorizontal_23_T & $signed(inSpriteXValue_23) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1040 = spriteScaleUpHorizontalReg_23 ? $signed({{2{_inSpriteX_23_T_4[10]}},_inSpriteX_23_T_4}) :
    $signed(_inSpriteX_23_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1041 = spriteScaleUpHorizontalReg_23 ? _inSpriteHorizontal_23_T_8 : _inSpriteHorizontal_23_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1042 = ~spriteScaleUpHorizontalReg_23 ? $signed({{1{inSpriteXValue_23[11]}},inSpriteXValue_23}) :
    $signed(_GEN_1040); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_23 = ~spriteScaleUpHorizontalReg_23 ? $signed(inSpriteXValue_23) >= 12'sh0 & $signed(
    inSpriteXValue_23) < 12'sh20 : _GEN_1041; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1797 = {{1{spriteYPositionReg_23[9]}},spriteYPositionReg_23}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_23 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1797); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_23 = inSpriteYValue_23[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_23_T = $signed(inSpriteYPreScaled_23) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_23_T_4 = inSpriteYPreScaled_23[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_23_T_8 = _inSpriteVertical_23_T & $signed(inSpriteYPreScaled_23) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_23_T_5 = {$signed(inSpriteYPreScaled_23), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_23_T_14 = _inSpriteVertical_23_T & $signed(inSpriteYPreScaled_23) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1048 = spriteScaleUpVerticalReg_23 ? $signed({{2{_inSpriteY_23_T_4[9]}},_inSpriteY_23_T_4}) :
    $signed(_inSpriteY_23_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1049 = spriteScaleUpVerticalReg_23 ? _inSpriteVertical_23_T_8 : _inSpriteVertical_23_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1050 = ~spriteScaleUpVerticalReg_23 ? $signed({{1{inSpriteYPreScaled_23[10]}},inSpriteYPreScaled_23})
     : $signed(_GEN_1048); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_23 = ~spriteScaleUpVerticalReg_23 ? $signed(inSpriteYPreScaled_23) >= 11'sh0 & $signed(
    inSpriteYPreScaled_23) < 11'sh20 : _GEN_1049; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_24 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_24); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_24_T = $signed(inSpriteXValue_24) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_24_T_4 = inSpriteXValue_24[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_24_T_8 = _inSpriteHorizontal_24_T & $signed(inSpriteXValue_24) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_24_T_5 = {$signed(inSpriteXValue_24), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_24_T_14 = _inSpriteHorizontal_24_T & $signed(inSpriteXValue_24) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1056 = spriteScaleUpHorizontalReg_24 ? $signed({{2{_inSpriteX_24_T_4[10]}},_inSpriteX_24_T_4}) :
    $signed(_inSpriteX_24_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1057 = spriteScaleUpHorizontalReg_24 ? _inSpriteHorizontal_24_T_8 : _inSpriteHorizontal_24_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1058 = ~spriteScaleUpHorizontalReg_24 ? $signed({{1{inSpriteXValue_24[11]}},inSpriteXValue_24}) :
    $signed(_GEN_1056); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_24 = ~spriteScaleUpHorizontalReg_24 ? $signed(inSpriteXValue_24) >= 12'sh0 & $signed(
    inSpriteXValue_24) < 12'sh20 : _GEN_1057; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1799 = {{1{spriteYPositionReg_24[9]}},spriteYPositionReg_24}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_24 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1799); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_24 = inSpriteYValue_24[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_24_T = $signed(inSpriteYPreScaled_24) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_24_T_4 = inSpriteYPreScaled_24[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_24_T_8 = _inSpriteVertical_24_T & $signed(inSpriteYPreScaled_24) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_24_T_5 = {$signed(inSpriteYPreScaled_24), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_24_T_14 = _inSpriteVertical_24_T & $signed(inSpriteYPreScaled_24) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1064 = spriteScaleUpVerticalReg_24 ? $signed({{2{_inSpriteY_24_T_4[9]}},_inSpriteY_24_T_4}) :
    $signed(_inSpriteY_24_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1065 = spriteScaleUpVerticalReg_24 ? _inSpriteVertical_24_T_8 : _inSpriteVertical_24_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1066 = ~spriteScaleUpVerticalReg_24 ? $signed({{1{inSpriteYPreScaled_24[10]}},inSpriteYPreScaled_24})
     : $signed(_GEN_1064); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_24 = ~spriteScaleUpVerticalReg_24 ? $signed(inSpriteYPreScaled_24) >= 11'sh0 & $signed(
    inSpriteYPreScaled_24) < 11'sh20 : _GEN_1065; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_25 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_25); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_25_T = $signed(inSpriteXValue_25) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_25_T_4 = inSpriteXValue_25[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_25_T_8 = _inSpriteHorizontal_25_T & $signed(inSpriteXValue_25) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_25_T_5 = {$signed(inSpriteXValue_25), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_25_T_14 = _inSpriteHorizontal_25_T & $signed(inSpriteXValue_25) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1072 = spriteScaleUpHorizontalReg_25 ? $signed({{2{_inSpriteX_25_T_4[10]}},_inSpriteX_25_T_4}) :
    $signed(_inSpriteX_25_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1073 = spriteScaleUpHorizontalReg_25 ? _inSpriteHorizontal_25_T_8 : _inSpriteHorizontal_25_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1074 = ~spriteScaleUpHorizontalReg_25 ? $signed({{1{inSpriteXValue_25[11]}},inSpriteXValue_25}) :
    $signed(_GEN_1072); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_25 = ~spriteScaleUpHorizontalReg_25 ? $signed(inSpriteXValue_25) >= 12'sh0 & $signed(
    inSpriteXValue_25) < 12'sh20 : _GEN_1073; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1801 = {{1{spriteYPositionReg_25[9]}},spriteYPositionReg_25}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_25 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1801); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_25 = inSpriteYValue_25[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_25_T = $signed(inSpriteYPreScaled_25) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_25_T_4 = inSpriteYPreScaled_25[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_25_T_8 = _inSpriteVertical_25_T & $signed(inSpriteYPreScaled_25) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_25_T_5 = {$signed(inSpriteYPreScaled_25), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_25_T_14 = _inSpriteVertical_25_T & $signed(inSpriteYPreScaled_25) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1080 = spriteScaleUpVerticalReg_25 ? $signed({{2{_inSpriteY_25_T_4[9]}},_inSpriteY_25_T_4}) :
    $signed(_inSpriteY_25_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1081 = spriteScaleUpVerticalReg_25 ? _inSpriteVertical_25_T_8 : _inSpriteVertical_25_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1082 = ~spriteScaleUpVerticalReg_25 ? $signed({{1{inSpriteYPreScaled_25[10]}},inSpriteYPreScaled_25})
     : $signed(_GEN_1080); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_25 = ~spriteScaleUpVerticalReg_25 ? $signed(inSpriteYPreScaled_25) >= 11'sh0 & $signed(
    inSpriteYPreScaled_25) < 11'sh20 : _GEN_1081; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_26 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_26); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_26_T = $signed(inSpriteXValue_26) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_26_T_4 = inSpriteXValue_26[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_26_T_8 = _inSpriteHorizontal_26_T & $signed(inSpriteXValue_26) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_26_T_5 = {$signed(inSpriteXValue_26), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_26_T_14 = _inSpriteHorizontal_26_T & $signed(inSpriteXValue_26) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1088 = spriteScaleUpHorizontalReg_26 ? $signed({{2{_inSpriteX_26_T_4[10]}},_inSpriteX_26_T_4}) :
    $signed(_inSpriteX_26_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1089 = spriteScaleUpHorizontalReg_26 ? _inSpriteHorizontal_26_T_8 : _inSpriteHorizontal_26_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1090 = ~spriteScaleUpHorizontalReg_26 ? $signed({{1{inSpriteXValue_26[11]}},inSpriteXValue_26}) :
    $signed(_GEN_1088); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_26 = ~spriteScaleUpHorizontalReg_26 ? $signed(inSpriteXValue_26) >= 12'sh0 & $signed(
    inSpriteXValue_26) < 12'sh20 : _GEN_1089; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1803 = {{1{spriteYPositionReg_26[9]}},spriteYPositionReg_26}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_26 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1803); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_26 = inSpriteYValue_26[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_26_T = $signed(inSpriteYPreScaled_26) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_26_T_4 = inSpriteYPreScaled_26[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_26_T_8 = _inSpriteVertical_26_T & $signed(inSpriteYPreScaled_26) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_26_T_5 = {$signed(inSpriteYPreScaled_26), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_26_T_14 = _inSpriteVertical_26_T & $signed(inSpriteYPreScaled_26) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1096 = spriteScaleUpVerticalReg_26 ? $signed({{2{_inSpriteY_26_T_4[9]}},_inSpriteY_26_T_4}) :
    $signed(_inSpriteY_26_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1097 = spriteScaleUpVerticalReg_26 ? _inSpriteVertical_26_T_8 : _inSpriteVertical_26_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1098 = ~spriteScaleUpVerticalReg_26 ? $signed({{1{inSpriteYPreScaled_26[10]}},inSpriteYPreScaled_26})
     : $signed(_GEN_1096); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_26 = ~spriteScaleUpVerticalReg_26 ? $signed(inSpriteYPreScaled_26) >= 11'sh0 & $signed(
    inSpriteYPreScaled_26) < 11'sh20 : _GEN_1097; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_27 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_27); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_27_T = $signed(inSpriteXValue_27) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_27_T_4 = inSpriteXValue_27[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_27_T_8 = _inSpriteHorizontal_27_T & $signed(inSpriteXValue_27) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_27_T_5 = {$signed(inSpriteXValue_27), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_27_T_14 = _inSpriteHorizontal_27_T & $signed(inSpriteXValue_27) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1104 = spriteScaleUpHorizontalReg_27 ? $signed({{2{_inSpriteX_27_T_4[10]}},_inSpriteX_27_T_4}) :
    $signed(_inSpriteX_27_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1105 = spriteScaleUpHorizontalReg_27 ? _inSpriteHorizontal_27_T_8 : _inSpriteHorizontal_27_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1106 = ~spriteScaleUpHorizontalReg_27 ? $signed({{1{inSpriteXValue_27[11]}},inSpriteXValue_27}) :
    $signed(_GEN_1104); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_27 = ~spriteScaleUpHorizontalReg_27 ? $signed(inSpriteXValue_27) >= 12'sh0 & $signed(
    inSpriteXValue_27) < 12'sh20 : _GEN_1105; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1805 = {{1{spriteYPositionReg_27[9]}},spriteYPositionReg_27}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_27 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1805); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_27 = inSpriteYValue_27[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_27_T = $signed(inSpriteYPreScaled_27) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_27_T_4 = inSpriteYPreScaled_27[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_27_T_8 = _inSpriteVertical_27_T & $signed(inSpriteYPreScaled_27) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_27_T_5 = {$signed(inSpriteYPreScaled_27), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_27_T_14 = _inSpriteVertical_27_T & $signed(inSpriteYPreScaled_27) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1112 = spriteScaleUpVerticalReg_27 ? $signed({{2{_inSpriteY_27_T_4[9]}},_inSpriteY_27_T_4}) :
    $signed(_inSpriteY_27_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1113 = spriteScaleUpVerticalReg_27 ? _inSpriteVertical_27_T_8 : _inSpriteVertical_27_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1114 = ~spriteScaleUpVerticalReg_27 ? $signed({{1{inSpriteYPreScaled_27[10]}},inSpriteYPreScaled_27})
     : $signed(_GEN_1112); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_27 = ~spriteScaleUpVerticalReg_27 ? $signed(inSpriteYPreScaled_27) >= 11'sh0 & $signed(
    inSpriteYPreScaled_27) < 11'sh20 : _GEN_1113; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_28 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_28); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_28_T = $signed(inSpriteXValue_28) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_28_T_4 = inSpriteXValue_28[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_28_T_8 = _inSpriteHorizontal_28_T & $signed(inSpriteXValue_28) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_28_T_5 = {$signed(inSpriteXValue_28), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_28_T_14 = _inSpriteHorizontal_28_T & $signed(inSpriteXValue_28) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1120 = spriteScaleUpHorizontalReg_28 ? $signed({{2{_inSpriteX_28_T_4[10]}},_inSpriteX_28_T_4}) :
    $signed(_inSpriteX_28_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1121 = spriteScaleUpHorizontalReg_28 ? _inSpriteHorizontal_28_T_8 : _inSpriteHorizontal_28_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1122 = ~spriteScaleUpHorizontalReg_28 ? $signed({{1{inSpriteXValue_28[11]}},inSpriteXValue_28}) :
    $signed(_GEN_1120); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_28 = ~spriteScaleUpHorizontalReg_28 ? $signed(inSpriteXValue_28) >= 12'sh0 & $signed(
    inSpriteXValue_28) < 12'sh20 : _GEN_1121; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1807 = {{1{spriteYPositionReg_28[9]}},spriteYPositionReg_28}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_28 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1807); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_28 = inSpriteYValue_28[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_28_T = $signed(inSpriteYPreScaled_28) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_28_T_4 = inSpriteYPreScaled_28[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_28_T_8 = _inSpriteVertical_28_T & $signed(inSpriteYPreScaled_28) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_28_T_5 = {$signed(inSpriteYPreScaled_28), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_28_T_14 = _inSpriteVertical_28_T & $signed(inSpriteYPreScaled_28) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1128 = spriteScaleUpVerticalReg_28 ? $signed({{2{_inSpriteY_28_T_4[9]}},_inSpriteY_28_T_4}) :
    $signed(_inSpriteY_28_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1129 = spriteScaleUpVerticalReg_28 ? _inSpriteVertical_28_T_8 : _inSpriteVertical_28_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1130 = ~spriteScaleUpVerticalReg_28 ? $signed({{1{inSpriteYPreScaled_28[10]}},inSpriteYPreScaled_28})
     : $signed(_GEN_1128); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_28 = ~spriteScaleUpVerticalReg_28 ? $signed(inSpriteYPreScaled_28) >= 11'sh0 & $signed(
    inSpriteYPreScaled_28) < 11'sh20 : _GEN_1129; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_29 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_29); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_29_T = $signed(inSpriteXValue_29) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_29_T_4 = inSpriteXValue_29[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_29_T_8 = _inSpriteHorizontal_29_T & $signed(inSpriteXValue_29) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_29_T_5 = {$signed(inSpriteXValue_29), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_29_T_14 = _inSpriteHorizontal_29_T & $signed(inSpriteXValue_29) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1136 = spriteScaleUpHorizontalReg_29 ? $signed({{2{_inSpriteX_29_T_4[10]}},_inSpriteX_29_T_4}) :
    $signed(_inSpriteX_29_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1137 = spriteScaleUpHorizontalReg_29 ? _inSpriteHorizontal_29_T_8 : _inSpriteHorizontal_29_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1138 = ~spriteScaleUpHorizontalReg_29 ? $signed({{1{inSpriteXValue_29[11]}},inSpriteXValue_29}) :
    $signed(_GEN_1136); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_29 = ~spriteScaleUpHorizontalReg_29 ? $signed(inSpriteXValue_29) >= 12'sh0 & $signed(
    inSpriteXValue_29) < 12'sh20 : _GEN_1137; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1809 = {{1{spriteYPositionReg_29[9]}},spriteYPositionReg_29}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_29 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1809); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_29 = inSpriteYValue_29[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_29_T = $signed(inSpriteYPreScaled_29) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_29_T_4 = inSpriteYPreScaled_29[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_29_T_8 = _inSpriteVertical_29_T & $signed(inSpriteYPreScaled_29) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_29_T_5 = {$signed(inSpriteYPreScaled_29), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_29_T_14 = _inSpriteVertical_29_T & $signed(inSpriteYPreScaled_29) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1144 = spriteScaleUpVerticalReg_29 ? $signed({{2{_inSpriteY_29_T_4[9]}},_inSpriteY_29_T_4}) :
    $signed(_inSpriteY_29_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1145 = spriteScaleUpVerticalReg_29 ? _inSpriteVertical_29_T_8 : _inSpriteVertical_29_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1146 = ~spriteScaleUpVerticalReg_29 ? $signed({{1{inSpriteYPreScaled_29[10]}},inSpriteYPreScaled_29})
     : $signed(_GEN_1144); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_29 = ~spriteScaleUpVerticalReg_29 ? $signed(inSpriteYPreScaled_29) >= 11'sh0 & $signed(
    inSpriteYPreScaled_29) < 11'sh20 : _GEN_1145; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_30 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_30); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_30_T = $signed(inSpriteXValue_30) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_30_T_4 = inSpriteXValue_30[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_30_T_8 = _inSpriteHorizontal_30_T & $signed(inSpriteXValue_30) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_30_T_5 = {$signed(inSpriteXValue_30), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_30_T_14 = _inSpriteHorizontal_30_T & $signed(inSpriteXValue_30) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1152 = spriteScaleUpHorizontalReg_30 ? $signed({{2{_inSpriteX_30_T_4[10]}},_inSpriteX_30_T_4}) :
    $signed(_inSpriteX_30_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1153 = spriteScaleUpHorizontalReg_30 ? _inSpriteHorizontal_30_T_8 : _inSpriteHorizontal_30_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1154 = ~spriteScaleUpHorizontalReg_30 ? $signed({{1{inSpriteXValue_30[11]}},inSpriteXValue_30}) :
    $signed(_GEN_1152); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_30 = ~spriteScaleUpHorizontalReg_30 ? $signed(inSpriteXValue_30) >= 12'sh0 & $signed(
    inSpriteXValue_30) < 12'sh20 : _GEN_1153; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1811 = {{1{spriteYPositionReg_30[9]}},spriteYPositionReg_30}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_30 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1811); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_30 = inSpriteYValue_30[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_30_T = $signed(inSpriteYPreScaled_30) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_30_T_4 = inSpriteYPreScaled_30[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_30_T_8 = _inSpriteVertical_30_T & $signed(inSpriteYPreScaled_30) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_30_T_5 = {$signed(inSpriteYPreScaled_30), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_30_T_14 = _inSpriteVertical_30_T & $signed(inSpriteYPreScaled_30) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1160 = spriteScaleUpVerticalReg_30 ? $signed({{2{_inSpriteY_30_T_4[9]}},_inSpriteY_30_T_4}) :
    $signed(_inSpriteY_30_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1161 = spriteScaleUpVerticalReg_30 ? _inSpriteVertical_30_T_8 : _inSpriteVertical_30_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1162 = ~spriteScaleUpVerticalReg_30 ? $signed({{1{inSpriteYPreScaled_30[10]}},inSpriteYPreScaled_30})
     : $signed(_GEN_1160); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_30 = ~spriteScaleUpVerticalReg_30 ? $signed(inSpriteYPreScaled_30) >= 11'sh0 & $signed(
    inSpriteYPreScaled_30) < 11'sh20 : _GEN_1161; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_31 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_31); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_31_T = $signed(inSpriteXValue_31) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_31_T_4 = inSpriteXValue_31[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_31_T_8 = _inSpriteHorizontal_31_T & $signed(inSpriteXValue_31) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_31_T_5 = {$signed(inSpriteXValue_31), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_31_T_14 = _inSpriteHorizontal_31_T & $signed(inSpriteXValue_31) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1168 = spriteScaleUpHorizontalReg_31 ? $signed({{2{_inSpriteX_31_T_4[10]}},_inSpriteX_31_T_4}) :
    $signed(_inSpriteX_31_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1169 = spriteScaleUpHorizontalReg_31 ? _inSpriteHorizontal_31_T_8 : _inSpriteHorizontal_31_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1170 = ~spriteScaleUpHorizontalReg_31 ? $signed({{1{inSpriteXValue_31[11]}},inSpriteXValue_31}) :
    $signed(_GEN_1168); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_31 = ~spriteScaleUpHorizontalReg_31 ? $signed(inSpriteXValue_31) >= 12'sh0 & $signed(
    inSpriteXValue_31) < 12'sh20 : _GEN_1169; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1813 = {{1{spriteYPositionReg_31[9]}},spriteYPositionReg_31}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_31 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1813); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_31 = inSpriteYValue_31[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_31_T = $signed(inSpriteYPreScaled_31) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_31_T_4 = inSpriteYPreScaled_31[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_31_T_8 = _inSpriteVertical_31_T & $signed(inSpriteYPreScaled_31) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_31_T_5 = {$signed(inSpriteYPreScaled_31), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_31_T_14 = _inSpriteVertical_31_T & $signed(inSpriteYPreScaled_31) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1176 = spriteScaleUpVerticalReg_31 ? $signed({{2{_inSpriteY_31_T_4[9]}},_inSpriteY_31_T_4}) :
    $signed(_inSpriteY_31_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1177 = spriteScaleUpVerticalReg_31 ? _inSpriteVertical_31_T_8 : _inSpriteVertical_31_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1178 = ~spriteScaleUpVerticalReg_31 ? $signed({{1{inSpriteYPreScaled_31[10]}},inSpriteYPreScaled_31})
     : $signed(_GEN_1176); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_31 = ~spriteScaleUpVerticalReg_31 ? $signed(inSpriteYPreScaled_31) >= 11'sh0 & $signed(
    inSpriteYPreScaled_31) < 11'sh20 : _GEN_1177; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_32 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_32); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_32_T = $signed(inSpriteXValue_32) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_32_T_4 = inSpriteXValue_32[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_32_T_8 = _inSpriteHorizontal_32_T & $signed(inSpriteXValue_32) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_32_T_5 = {$signed(inSpriteXValue_32), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_32_T_14 = _inSpriteHorizontal_32_T & $signed(inSpriteXValue_32) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1184 = spriteScaleUpHorizontalReg_32 ? $signed({{2{_inSpriteX_32_T_4[10]}},_inSpriteX_32_T_4}) :
    $signed(_inSpriteX_32_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1185 = spriteScaleUpHorizontalReg_32 ? _inSpriteHorizontal_32_T_8 : _inSpriteHorizontal_32_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1186 = ~spriteScaleUpHorizontalReg_32 ? $signed({{1{inSpriteXValue_32[11]}},inSpriteXValue_32}) :
    $signed(_GEN_1184); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_32 = ~spriteScaleUpHorizontalReg_32 ? $signed(inSpriteXValue_32) >= 12'sh0 & $signed(
    inSpriteXValue_32) < 12'sh20 : _GEN_1185; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1815 = {{1{spriteYPositionReg_32[9]}},spriteYPositionReg_32}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_32 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1815); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_32 = inSpriteYValue_32[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_32_T = $signed(inSpriteYPreScaled_32) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_32_T_4 = inSpriteYPreScaled_32[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_32_T_8 = _inSpriteVertical_32_T & $signed(inSpriteYPreScaled_32) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_32_T_5 = {$signed(inSpriteYPreScaled_32), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_32_T_14 = _inSpriteVertical_32_T & $signed(inSpriteYPreScaled_32) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1192 = spriteScaleUpVerticalReg_32 ? $signed({{2{_inSpriteY_32_T_4[9]}},_inSpriteY_32_T_4}) :
    $signed(_inSpriteY_32_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1193 = spriteScaleUpVerticalReg_32 ? _inSpriteVertical_32_T_8 : _inSpriteVertical_32_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1194 = ~spriteScaleUpVerticalReg_32 ? $signed({{1{inSpriteYPreScaled_32[10]}},inSpriteYPreScaled_32})
     : $signed(_GEN_1192); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_32 = ~spriteScaleUpVerticalReg_32 ? $signed(inSpriteYPreScaled_32) >= 11'sh0 & $signed(
    inSpriteYPreScaled_32) < 11'sh20 : _GEN_1193; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_33 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_33); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_33_T = $signed(inSpriteXValue_33) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_33_T_4 = inSpriteXValue_33[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_33_T_8 = _inSpriteHorizontal_33_T & $signed(inSpriteXValue_33) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_33_T_5 = {$signed(inSpriteXValue_33), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_33_T_14 = _inSpriteHorizontal_33_T & $signed(inSpriteXValue_33) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1200 = spriteScaleUpHorizontalReg_33 ? $signed({{2{_inSpriteX_33_T_4[10]}},_inSpriteX_33_T_4}) :
    $signed(_inSpriteX_33_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1201 = spriteScaleUpHorizontalReg_33 ? _inSpriteHorizontal_33_T_8 : _inSpriteHorizontal_33_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1202 = ~spriteScaleUpHorizontalReg_33 ? $signed({{1{inSpriteXValue_33[11]}},inSpriteXValue_33}) :
    $signed(_GEN_1200); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_33 = ~spriteScaleUpHorizontalReg_33 ? $signed(inSpriteXValue_33) >= 12'sh0 & $signed(
    inSpriteXValue_33) < 12'sh20 : _GEN_1201; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1817 = {{1{spriteYPositionReg_33[9]}},spriteYPositionReg_33}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_33 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1817); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_33 = inSpriteYValue_33[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_33_T = $signed(inSpriteYPreScaled_33) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_33_T_4 = inSpriteYPreScaled_33[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_33_T_8 = _inSpriteVertical_33_T & $signed(inSpriteYPreScaled_33) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_33_T_5 = {$signed(inSpriteYPreScaled_33), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_33_T_14 = _inSpriteVertical_33_T & $signed(inSpriteYPreScaled_33) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1208 = spriteScaleUpVerticalReg_33 ? $signed({{2{_inSpriteY_33_T_4[9]}},_inSpriteY_33_T_4}) :
    $signed(_inSpriteY_33_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1209 = spriteScaleUpVerticalReg_33 ? _inSpriteVertical_33_T_8 : _inSpriteVertical_33_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1210 = ~spriteScaleUpVerticalReg_33 ? $signed({{1{inSpriteYPreScaled_33[10]}},inSpriteYPreScaled_33})
     : $signed(_GEN_1208); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_33 = ~spriteScaleUpVerticalReg_33 ? $signed(inSpriteYPreScaled_33) >= 11'sh0 & $signed(
    inSpriteYPreScaled_33) < 11'sh20 : _GEN_1209; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_34 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_34); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_34_T = $signed(inSpriteXValue_34) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_34_T_4 = inSpriteXValue_34[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_34_T_8 = _inSpriteHorizontal_34_T & $signed(inSpriteXValue_34) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_34_T_5 = {$signed(inSpriteXValue_34), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_34_T_14 = _inSpriteHorizontal_34_T & $signed(inSpriteXValue_34) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1216 = spriteScaleUpHorizontalReg_34 ? $signed({{2{_inSpriteX_34_T_4[10]}},_inSpriteX_34_T_4}) :
    $signed(_inSpriteX_34_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1217 = spriteScaleUpHorizontalReg_34 ? _inSpriteHorizontal_34_T_8 : _inSpriteHorizontal_34_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1218 = ~spriteScaleUpHorizontalReg_34 ? $signed({{1{inSpriteXValue_34[11]}},inSpriteXValue_34}) :
    $signed(_GEN_1216); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_34 = ~spriteScaleUpHorizontalReg_34 ? $signed(inSpriteXValue_34) >= 12'sh0 & $signed(
    inSpriteXValue_34) < 12'sh20 : _GEN_1217; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1819 = {{1{spriteYPositionReg_34[9]}},spriteYPositionReg_34}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_34 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1819); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_34 = inSpriteYValue_34[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_34_T = $signed(inSpriteYPreScaled_34) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_34_T_4 = inSpriteYPreScaled_34[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_34_T_8 = _inSpriteVertical_34_T & $signed(inSpriteYPreScaled_34) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_34_T_5 = {$signed(inSpriteYPreScaled_34), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_34_T_14 = _inSpriteVertical_34_T & $signed(inSpriteYPreScaled_34) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1224 = spriteScaleUpVerticalReg_34 ? $signed({{2{_inSpriteY_34_T_4[9]}},_inSpriteY_34_T_4}) :
    $signed(_inSpriteY_34_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1225 = spriteScaleUpVerticalReg_34 ? _inSpriteVertical_34_T_8 : _inSpriteVertical_34_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1226 = ~spriteScaleUpVerticalReg_34 ? $signed({{1{inSpriteYPreScaled_34[10]}},inSpriteYPreScaled_34})
     : $signed(_GEN_1224); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_34 = ~spriteScaleUpVerticalReg_34 ? $signed(inSpriteYPreScaled_34) >= 11'sh0 & $signed(
    inSpriteYPreScaled_34) < 11'sh20 : _GEN_1225; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_35 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_35); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_35_T = $signed(inSpriteXValue_35) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_35_T_4 = inSpriteXValue_35[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_35_T_8 = _inSpriteHorizontal_35_T & $signed(inSpriteXValue_35) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_35_T_5 = {$signed(inSpriteXValue_35), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_35_T_14 = _inSpriteHorizontal_35_T & $signed(inSpriteXValue_35) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1232 = spriteScaleUpHorizontalReg_35 ? $signed({{2{_inSpriteX_35_T_4[10]}},_inSpriteX_35_T_4}) :
    $signed(_inSpriteX_35_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1233 = spriteScaleUpHorizontalReg_35 ? _inSpriteHorizontal_35_T_8 : _inSpriteHorizontal_35_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1234 = ~spriteScaleUpHorizontalReg_35 ? $signed({{1{inSpriteXValue_35[11]}},inSpriteXValue_35}) :
    $signed(_GEN_1232); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_35 = ~spriteScaleUpHorizontalReg_35 ? $signed(inSpriteXValue_35) >= 12'sh0 & $signed(
    inSpriteXValue_35) < 12'sh20 : _GEN_1233; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1821 = {{1{spriteYPositionReg_35[9]}},spriteYPositionReg_35}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_35 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1821); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_35 = inSpriteYValue_35[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_35_T = $signed(inSpriteYPreScaled_35) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_35_T_4 = inSpriteYPreScaled_35[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_35_T_8 = _inSpriteVertical_35_T & $signed(inSpriteYPreScaled_35) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_35_T_5 = {$signed(inSpriteYPreScaled_35), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_35_T_14 = _inSpriteVertical_35_T & $signed(inSpriteYPreScaled_35) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1240 = spriteScaleUpVerticalReg_35 ? $signed({{2{_inSpriteY_35_T_4[9]}},_inSpriteY_35_T_4}) :
    $signed(_inSpriteY_35_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1241 = spriteScaleUpVerticalReg_35 ? _inSpriteVertical_35_T_8 : _inSpriteVertical_35_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1242 = ~spriteScaleUpVerticalReg_35 ? $signed({{1{inSpriteYPreScaled_35[10]}},inSpriteYPreScaled_35})
     : $signed(_GEN_1240); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_35 = ~spriteScaleUpVerticalReg_35 ? $signed(inSpriteYPreScaled_35) >= 11'sh0 & $signed(
    inSpriteYPreScaled_35) < 11'sh20 : _GEN_1241; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_36 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_36); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_36_T = $signed(inSpriteXValue_36) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_36_T_4 = inSpriteXValue_36[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_36_T_8 = _inSpriteHorizontal_36_T & $signed(inSpriteXValue_36) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_36_T_5 = {$signed(inSpriteXValue_36), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_36_T_14 = _inSpriteHorizontal_36_T & $signed(inSpriteXValue_36) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1248 = spriteScaleUpHorizontalReg_36 ? $signed({{2{_inSpriteX_36_T_4[10]}},_inSpriteX_36_T_4}) :
    $signed(_inSpriteX_36_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1249 = spriteScaleUpHorizontalReg_36 ? _inSpriteHorizontal_36_T_8 : _inSpriteHorizontal_36_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1250 = ~spriteScaleUpHorizontalReg_36 ? $signed({{1{inSpriteXValue_36[11]}},inSpriteXValue_36}) :
    $signed(_GEN_1248); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_36 = ~spriteScaleUpHorizontalReg_36 ? $signed(inSpriteXValue_36) >= 12'sh0 & $signed(
    inSpriteXValue_36) < 12'sh20 : _GEN_1249; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1823 = {{1{spriteYPositionReg_36[9]}},spriteYPositionReg_36}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_36 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1823); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_36 = inSpriteYValue_36[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_36_T = $signed(inSpriteYPreScaled_36) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_36_T_4 = inSpriteYPreScaled_36[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_36_T_8 = _inSpriteVertical_36_T & $signed(inSpriteYPreScaled_36) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_36_T_5 = {$signed(inSpriteYPreScaled_36), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_36_T_14 = _inSpriteVertical_36_T & $signed(inSpriteYPreScaled_36) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1256 = spriteScaleUpVerticalReg_36 ? $signed({{2{_inSpriteY_36_T_4[9]}},_inSpriteY_36_T_4}) :
    $signed(_inSpriteY_36_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1257 = spriteScaleUpVerticalReg_36 ? _inSpriteVertical_36_T_8 : _inSpriteVertical_36_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1258 = ~spriteScaleUpVerticalReg_36 ? $signed({{1{inSpriteYPreScaled_36[10]}},inSpriteYPreScaled_36})
     : $signed(_GEN_1256); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_36 = ~spriteScaleUpVerticalReg_36 ? $signed(inSpriteYPreScaled_36) >= 11'sh0 & $signed(
    inSpriteYPreScaled_36) < 11'sh20 : _GEN_1257; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_37 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_37); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_37_T = $signed(inSpriteXValue_37) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_37_T_4 = inSpriteXValue_37[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_37_T_8 = _inSpriteHorizontal_37_T & $signed(inSpriteXValue_37) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_37_T_5 = {$signed(inSpriteXValue_37), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_37_T_14 = _inSpriteHorizontal_37_T & $signed(inSpriteXValue_37) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1264 = spriteScaleUpHorizontalReg_37 ? $signed({{2{_inSpriteX_37_T_4[10]}},_inSpriteX_37_T_4}) :
    $signed(_inSpriteX_37_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1265 = spriteScaleUpHorizontalReg_37 ? _inSpriteHorizontal_37_T_8 : _inSpriteHorizontal_37_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1266 = ~spriteScaleUpHorizontalReg_37 ? $signed({{1{inSpriteXValue_37[11]}},inSpriteXValue_37}) :
    $signed(_GEN_1264); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_37 = ~spriteScaleUpHorizontalReg_37 ? $signed(inSpriteXValue_37) >= 12'sh0 & $signed(
    inSpriteXValue_37) < 12'sh20 : _GEN_1265; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1825 = {{1{spriteYPositionReg_37[9]}},spriteYPositionReg_37}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_37 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1825); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_37 = inSpriteYValue_37[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_37_T = $signed(inSpriteYPreScaled_37) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_37_T_4 = inSpriteYPreScaled_37[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_37_T_8 = _inSpriteVertical_37_T & $signed(inSpriteYPreScaled_37) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_37_T_5 = {$signed(inSpriteYPreScaled_37), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_37_T_14 = _inSpriteVertical_37_T & $signed(inSpriteYPreScaled_37) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1272 = spriteScaleUpVerticalReg_37 ? $signed({{2{_inSpriteY_37_T_4[9]}},_inSpriteY_37_T_4}) :
    $signed(_inSpriteY_37_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1273 = spriteScaleUpVerticalReg_37 ? _inSpriteVertical_37_T_8 : _inSpriteVertical_37_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1274 = ~spriteScaleUpVerticalReg_37 ? $signed({{1{inSpriteYPreScaled_37[10]}},inSpriteYPreScaled_37})
     : $signed(_GEN_1272); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_37 = ~spriteScaleUpVerticalReg_37 ? $signed(inSpriteYPreScaled_37) >= 11'sh0 & $signed(
    inSpriteYPreScaled_37) < 11'sh20 : _GEN_1273; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_38 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_38); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_38_T = $signed(inSpriteXValue_38) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_38_T_4 = inSpriteXValue_38[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_38_T_8 = _inSpriteHorizontal_38_T & $signed(inSpriteXValue_38) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_38_T_5 = {$signed(inSpriteXValue_38), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_38_T_14 = _inSpriteHorizontal_38_T & $signed(inSpriteXValue_38) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1280 = spriteScaleUpHorizontalReg_38 ? $signed({{2{_inSpriteX_38_T_4[10]}},_inSpriteX_38_T_4}) :
    $signed(_inSpriteX_38_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1281 = spriteScaleUpHorizontalReg_38 ? _inSpriteHorizontal_38_T_8 : _inSpriteHorizontal_38_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1282 = ~spriteScaleUpHorizontalReg_38 ? $signed({{1{inSpriteXValue_38[11]}},inSpriteXValue_38}) :
    $signed(_GEN_1280); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_38 = ~spriteScaleUpHorizontalReg_38 ? $signed(inSpriteXValue_38) >= 12'sh0 & $signed(
    inSpriteXValue_38) < 12'sh20 : _GEN_1281; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1827 = {{1{spriteYPositionReg_38[9]}},spriteYPositionReg_38}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_38 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1827); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_38 = inSpriteYValue_38[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_38_T = $signed(inSpriteYPreScaled_38) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_38_T_4 = inSpriteYPreScaled_38[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_38_T_8 = _inSpriteVertical_38_T & $signed(inSpriteYPreScaled_38) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_38_T_5 = {$signed(inSpriteYPreScaled_38), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_38_T_14 = _inSpriteVertical_38_T & $signed(inSpriteYPreScaled_38) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1288 = spriteScaleUpVerticalReg_38 ? $signed({{2{_inSpriteY_38_T_4[9]}},_inSpriteY_38_T_4}) :
    $signed(_inSpriteY_38_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1289 = spriteScaleUpVerticalReg_38 ? _inSpriteVertical_38_T_8 : _inSpriteVertical_38_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1290 = ~spriteScaleUpVerticalReg_38 ? $signed({{1{inSpriteYPreScaled_38[10]}},inSpriteYPreScaled_38})
     : $signed(_GEN_1288); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_38 = ~spriteScaleUpVerticalReg_38 ? $signed(inSpriteYPreScaled_38) >= 11'sh0 & $signed(
    inSpriteYPreScaled_38) < 11'sh20 : _GEN_1289; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_39 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_39); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_39_T = $signed(inSpriteXValue_39) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_39_T_4 = inSpriteXValue_39[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_39_T_8 = _inSpriteHorizontal_39_T & $signed(inSpriteXValue_39) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_39_T_5 = {$signed(inSpriteXValue_39), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_39_T_14 = _inSpriteHorizontal_39_T & $signed(inSpriteXValue_39) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1296 = spriteScaleUpHorizontalReg_39 ? $signed({{2{_inSpriteX_39_T_4[10]}},_inSpriteX_39_T_4}) :
    $signed(_inSpriteX_39_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1297 = spriteScaleUpHorizontalReg_39 ? _inSpriteHorizontal_39_T_8 : _inSpriteHorizontal_39_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1298 = ~spriteScaleUpHorizontalReg_39 ? $signed({{1{inSpriteXValue_39[11]}},inSpriteXValue_39}) :
    $signed(_GEN_1296); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_39 = ~spriteScaleUpHorizontalReg_39 ? $signed(inSpriteXValue_39) >= 12'sh0 & $signed(
    inSpriteXValue_39) < 12'sh20 : _GEN_1297; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1829 = {{1{spriteYPositionReg_39[9]}},spriteYPositionReg_39}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_39 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1829); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_39 = inSpriteYValue_39[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_39_T = $signed(inSpriteYPreScaled_39) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_39_T_4 = inSpriteYPreScaled_39[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_39_T_8 = _inSpriteVertical_39_T & $signed(inSpriteYPreScaled_39) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_39_T_5 = {$signed(inSpriteYPreScaled_39), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_39_T_14 = _inSpriteVertical_39_T & $signed(inSpriteYPreScaled_39) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1304 = spriteScaleUpVerticalReg_39 ? $signed({{2{_inSpriteY_39_T_4[9]}},_inSpriteY_39_T_4}) :
    $signed(_inSpriteY_39_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1305 = spriteScaleUpVerticalReg_39 ? _inSpriteVertical_39_T_8 : _inSpriteVertical_39_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1306 = ~spriteScaleUpVerticalReg_39 ? $signed({{1{inSpriteYPreScaled_39[10]}},inSpriteYPreScaled_39})
     : $signed(_GEN_1304); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_39 = ~spriteScaleUpVerticalReg_39 ? $signed(inSpriteYPreScaled_39) >= 11'sh0 & $signed(
    inSpriteYPreScaled_39) < 11'sh20 : _GEN_1305; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_40 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_40); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_40_T = $signed(inSpriteXValue_40) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_40_T_4 = inSpriteXValue_40[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_40_T_8 = _inSpriteHorizontal_40_T & $signed(inSpriteXValue_40) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_40_T_5 = {$signed(inSpriteXValue_40), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_40_T_14 = _inSpriteHorizontal_40_T & $signed(inSpriteXValue_40) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1312 = spriteScaleUpHorizontalReg_40 ? $signed({{2{_inSpriteX_40_T_4[10]}},_inSpriteX_40_T_4}) :
    $signed(_inSpriteX_40_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1313 = spriteScaleUpHorizontalReg_40 ? _inSpriteHorizontal_40_T_8 : _inSpriteHorizontal_40_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1314 = ~spriteScaleUpHorizontalReg_40 ? $signed({{1{inSpriteXValue_40[11]}},inSpriteXValue_40}) :
    $signed(_GEN_1312); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_40 = ~spriteScaleUpHorizontalReg_40 ? $signed(inSpriteXValue_40) >= 12'sh0 & $signed(
    inSpriteXValue_40) < 12'sh20 : _GEN_1313; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1831 = {{1{spriteYPositionReg_40[9]}},spriteYPositionReg_40}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_40 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1831); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_40 = inSpriteYValue_40[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_40_T = $signed(inSpriteYPreScaled_40) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_40_T_4 = inSpriteYPreScaled_40[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_40_T_8 = _inSpriteVertical_40_T & $signed(inSpriteYPreScaled_40) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_40_T_5 = {$signed(inSpriteYPreScaled_40), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_40_T_14 = _inSpriteVertical_40_T & $signed(inSpriteYPreScaled_40) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1320 = spriteScaleUpVerticalReg_40 ? $signed({{2{_inSpriteY_40_T_4[9]}},_inSpriteY_40_T_4}) :
    $signed(_inSpriteY_40_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1321 = spriteScaleUpVerticalReg_40 ? _inSpriteVertical_40_T_8 : _inSpriteVertical_40_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1322 = ~spriteScaleUpVerticalReg_40 ? $signed({{1{inSpriteYPreScaled_40[10]}},inSpriteYPreScaled_40})
     : $signed(_GEN_1320); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_40 = ~spriteScaleUpVerticalReg_40 ? $signed(inSpriteYPreScaled_40) >= 11'sh0 & $signed(
    inSpriteYPreScaled_40) < 11'sh20 : _GEN_1321; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_41 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_41); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_41_T = $signed(inSpriteXValue_41) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_41_T_4 = inSpriteXValue_41[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_41_T_8 = _inSpriteHorizontal_41_T & $signed(inSpriteXValue_41) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_41_T_5 = {$signed(inSpriteXValue_41), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_41_T_14 = _inSpriteHorizontal_41_T & $signed(inSpriteXValue_41) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1328 = spriteScaleUpHorizontalReg_41 ? $signed({{2{_inSpriteX_41_T_4[10]}},_inSpriteX_41_T_4}) :
    $signed(_inSpriteX_41_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1329 = spriteScaleUpHorizontalReg_41 ? _inSpriteHorizontal_41_T_8 : _inSpriteHorizontal_41_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1330 = ~spriteScaleUpHorizontalReg_41 ? $signed({{1{inSpriteXValue_41[11]}},inSpriteXValue_41}) :
    $signed(_GEN_1328); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_41 = ~spriteScaleUpHorizontalReg_41 ? $signed(inSpriteXValue_41) >= 12'sh0 & $signed(
    inSpriteXValue_41) < 12'sh20 : _GEN_1329; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1833 = {{1{spriteYPositionReg_41[9]}},spriteYPositionReg_41}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_41 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1833); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_41 = inSpriteYValue_41[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_41_T = $signed(inSpriteYPreScaled_41) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_41_T_4 = inSpriteYPreScaled_41[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_41_T_8 = _inSpriteVertical_41_T & $signed(inSpriteYPreScaled_41) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_41_T_5 = {$signed(inSpriteYPreScaled_41), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_41_T_14 = _inSpriteVertical_41_T & $signed(inSpriteYPreScaled_41) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1336 = spriteScaleUpVerticalReg_41 ? $signed({{2{_inSpriteY_41_T_4[9]}},_inSpriteY_41_T_4}) :
    $signed(_inSpriteY_41_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1337 = spriteScaleUpVerticalReg_41 ? _inSpriteVertical_41_T_8 : _inSpriteVertical_41_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1338 = ~spriteScaleUpVerticalReg_41 ? $signed({{1{inSpriteYPreScaled_41[10]}},inSpriteYPreScaled_41})
     : $signed(_GEN_1336); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_41 = ~spriteScaleUpVerticalReg_41 ? $signed(inSpriteYPreScaled_41) >= 11'sh0 & $signed(
    inSpriteYPreScaled_41) < 11'sh20 : _GEN_1337; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_42 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_42); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_42_T = $signed(inSpriteXValue_42) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_42_T_4 = inSpriteXValue_42[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_42_T_8 = _inSpriteHorizontal_42_T & $signed(inSpriteXValue_42) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_42_T_5 = {$signed(inSpriteXValue_42), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_42_T_14 = _inSpriteHorizontal_42_T & $signed(inSpriteXValue_42) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1344 = spriteScaleUpHorizontalReg_42 ? $signed({{2{_inSpriteX_42_T_4[10]}},_inSpriteX_42_T_4}) :
    $signed(_inSpriteX_42_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1345 = spriteScaleUpHorizontalReg_42 ? _inSpriteHorizontal_42_T_8 : _inSpriteHorizontal_42_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1346 = ~spriteScaleUpHorizontalReg_42 ? $signed({{1{inSpriteXValue_42[11]}},inSpriteXValue_42}) :
    $signed(_GEN_1344); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_42 = ~spriteScaleUpHorizontalReg_42 ? $signed(inSpriteXValue_42) >= 12'sh0 & $signed(
    inSpriteXValue_42) < 12'sh20 : _GEN_1345; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1835 = {{1{spriteYPositionReg_42[9]}},spriteYPositionReg_42}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_42 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1835); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_42 = inSpriteYValue_42[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_42_T = $signed(inSpriteYPreScaled_42) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_42_T_4 = inSpriteYPreScaled_42[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_42_T_8 = _inSpriteVertical_42_T & $signed(inSpriteYPreScaled_42) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_42_T_5 = {$signed(inSpriteYPreScaled_42), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_42_T_14 = _inSpriteVertical_42_T & $signed(inSpriteYPreScaled_42) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1352 = spriteScaleUpVerticalReg_42 ? $signed({{2{_inSpriteY_42_T_4[9]}},_inSpriteY_42_T_4}) :
    $signed(_inSpriteY_42_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1353 = spriteScaleUpVerticalReg_42 ? _inSpriteVertical_42_T_8 : _inSpriteVertical_42_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1354 = ~spriteScaleUpVerticalReg_42 ? $signed({{1{inSpriteYPreScaled_42[10]}},inSpriteYPreScaled_42})
     : $signed(_GEN_1352); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_42 = ~spriteScaleUpVerticalReg_42 ? $signed(inSpriteYPreScaled_42) >= 11'sh0 & $signed(
    inSpriteYPreScaled_42) < 11'sh20 : _GEN_1353; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_43 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_43); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_43_T = $signed(inSpriteXValue_43) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_43_T_4 = inSpriteXValue_43[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_43_T_8 = _inSpriteHorizontal_43_T & $signed(inSpriteXValue_43) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_43_T_5 = {$signed(inSpriteXValue_43), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_43_T_14 = _inSpriteHorizontal_43_T & $signed(inSpriteXValue_43) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1360 = spriteScaleUpHorizontalReg_43 ? $signed({{2{_inSpriteX_43_T_4[10]}},_inSpriteX_43_T_4}) :
    $signed(_inSpriteX_43_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1361 = spriteScaleUpHorizontalReg_43 ? _inSpriteHorizontal_43_T_8 : _inSpriteHorizontal_43_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1362 = ~spriteScaleUpHorizontalReg_43 ? $signed({{1{inSpriteXValue_43[11]}},inSpriteXValue_43}) :
    $signed(_GEN_1360); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_43 = ~spriteScaleUpHorizontalReg_43 ? $signed(inSpriteXValue_43) >= 12'sh0 & $signed(
    inSpriteXValue_43) < 12'sh20 : _GEN_1361; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1837 = {{1{spriteYPositionReg_43[9]}},spriteYPositionReg_43}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_43 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1837); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_43 = inSpriteYValue_43[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_43_T = $signed(inSpriteYPreScaled_43) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_43_T_4 = inSpriteYPreScaled_43[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_43_T_8 = _inSpriteVertical_43_T & $signed(inSpriteYPreScaled_43) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_43_T_5 = {$signed(inSpriteYPreScaled_43), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_43_T_14 = _inSpriteVertical_43_T & $signed(inSpriteYPreScaled_43) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1368 = spriteScaleUpVerticalReg_43 ? $signed({{2{_inSpriteY_43_T_4[9]}},_inSpriteY_43_T_4}) :
    $signed(_inSpriteY_43_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1369 = spriteScaleUpVerticalReg_43 ? _inSpriteVertical_43_T_8 : _inSpriteVertical_43_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1370 = ~spriteScaleUpVerticalReg_43 ? $signed({{1{inSpriteYPreScaled_43[10]}},inSpriteYPreScaled_43})
     : $signed(_GEN_1368); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_43 = ~spriteScaleUpVerticalReg_43 ? $signed(inSpriteYPreScaled_43) >= 11'sh0 & $signed(
    inSpriteYPreScaled_43) < 11'sh20 : _GEN_1369; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_44 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_44); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_44_T = $signed(inSpriteXValue_44) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_44_T_4 = inSpriteXValue_44[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_44_T_8 = _inSpriteHorizontal_44_T & $signed(inSpriteXValue_44) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_44_T_5 = {$signed(inSpriteXValue_44), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_44_T_14 = _inSpriteHorizontal_44_T & $signed(inSpriteXValue_44) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1376 = spriteScaleUpHorizontalReg_44 ? $signed({{2{_inSpriteX_44_T_4[10]}},_inSpriteX_44_T_4}) :
    $signed(_inSpriteX_44_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1377 = spriteScaleUpHorizontalReg_44 ? _inSpriteHorizontal_44_T_8 : _inSpriteHorizontal_44_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1378 = ~spriteScaleUpHorizontalReg_44 ? $signed({{1{inSpriteXValue_44[11]}},inSpriteXValue_44}) :
    $signed(_GEN_1376); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_44 = ~spriteScaleUpHorizontalReg_44 ? $signed(inSpriteXValue_44) >= 12'sh0 & $signed(
    inSpriteXValue_44) < 12'sh20 : _GEN_1377; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1839 = {{1{spriteYPositionReg_44[9]}},spriteYPositionReg_44}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_44 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1839); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_44 = inSpriteYValue_44[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_44_T = $signed(inSpriteYPreScaled_44) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_44_T_4 = inSpriteYPreScaled_44[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_44_T_8 = _inSpriteVertical_44_T & $signed(inSpriteYPreScaled_44) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_44_T_5 = {$signed(inSpriteYPreScaled_44), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_44_T_14 = _inSpriteVertical_44_T & $signed(inSpriteYPreScaled_44) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1384 = spriteScaleUpVerticalReg_44 ? $signed({{2{_inSpriteY_44_T_4[9]}},_inSpriteY_44_T_4}) :
    $signed(_inSpriteY_44_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1385 = spriteScaleUpVerticalReg_44 ? _inSpriteVertical_44_T_8 : _inSpriteVertical_44_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1386 = ~spriteScaleUpVerticalReg_44 ? $signed({{1{inSpriteYPreScaled_44[10]}},inSpriteYPreScaled_44})
     : $signed(_GEN_1384); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_44 = ~spriteScaleUpVerticalReg_44 ? $signed(inSpriteYPreScaled_44) >= 11'sh0 & $signed(
    inSpriteYPreScaled_44) < 11'sh20 : _GEN_1385; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_45 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_45); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_45_T = $signed(inSpriteXValue_45) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_45_T_4 = inSpriteXValue_45[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_45_T_8 = _inSpriteHorizontal_45_T & $signed(inSpriteXValue_45) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_45_T_5 = {$signed(inSpriteXValue_45), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_45_T_14 = _inSpriteHorizontal_45_T & $signed(inSpriteXValue_45) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1392 = spriteScaleUpHorizontalReg_45 ? $signed({{2{_inSpriteX_45_T_4[10]}},_inSpriteX_45_T_4}) :
    $signed(_inSpriteX_45_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1393 = spriteScaleUpHorizontalReg_45 ? _inSpriteHorizontal_45_T_8 : _inSpriteHorizontal_45_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1394 = ~spriteScaleUpHorizontalReg_45 ? $signed({{1{inSpriteXValue_45[11]}},inSpriteXValue_45}) :
    $signed(_GEN_1392); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_45 = ~spriteScaleUpHorizontalReg_45 ? $signed(inSpriteXValue_45) >= 12'sh0 & $signed(
    inSpriteXValue_45) < 12'sh20 : _GEN_1393; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1841 = {{1{spriteYPositionReg_45[9]}},spriteYPositionReg_45}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_45 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1841); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_45 = inSpriteYValue_45[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_45_T = $signed(inSpriteYPreScaled_45) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_45_T_4 = inSpriteYPreScaled_45[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_45_T_8 = _inSpriteVertical_45_T & $signed(inSpriteYPreScaled_45) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_45_T_5 = {$signed(inSpriteYPreScaled_45), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_45_T_14 = _inSpriteVertical_45_T & $signed(inSpriteYPreScaled_45) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1400 = spriteScaleUpVerticalReg_45 ? $signed({{2{_inSpriteY_45_T_4[9]}},_inSpriteY_45_T_4}) :
    $signed(_inSpriteY_45_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1401 = spriteScaleUpVerticalReg_45 ? _inSpriteVertical_45_T_8 : _inSpriteVertical_45_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1402 = ~spriteScaleUpVerticalReg_45 ? $signed({{1{inSpriteYPreScaled_45[10]}},inSpriteYPreScaled_45})
     : $signed(_GEN_1400); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_45 = ~spriteScaleUpVerticalReg_45 ? $signed(inSpriteYPreScaled_45) >= 11'sh0 & $signed(
    inSpriteYPreScaled_45) < 11'sh20 : _GEN_1401; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_46 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_46); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_46 = $signed(inSpriteXValue_46) >= 12'sh0 & $signed(inSpriteXValue_46) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1410 = {{1{inSpriteXValue_46[11]}},inSpriteXValue_46}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1843 = {{1{spriteYPositionReg_46[9]}},spriteYPositionReg_46}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_46 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1843); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_46 = inSpriteYValue_46[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_46 = $signed(inSpriteYPreScaled_46) >= 11'sh0 & $signed(inSpriteYPreScaled_46) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1418 = {{1{inSpriteYPreScaled_46[10]}},inSpriteYPreScaled_46}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_47 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_47); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_47 = $signed(inSpriteXValue_47) >= 12'sh0 & $signed(inSpriteXValue_47) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1426 = {{1{inSpriteXValue_47[11]}},inSpriteXValue_47}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1845 = {{1{spriteYPositionReg_47[9]}},spriteYPositionReg_47}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_47 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1845); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_47 = inSpriteYValue_47[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_47 = $signed(inSpriteYPreScaled_47) >= 11'sh0 & $signed(inSpriteYPreScaled_47) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1434 = {{1{inSpriteYPreScaled_47[10]}},inSpriteYPreScaled_47}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_48 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_48); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_48 = $signed(inSpriteXValue_48) >= 12'sh0 & $signed(inSpriteXValue_48) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1442 = {{1{inSpriteXValue_48[11]}},inSpriteXValue_48}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1847 = {{1{spriteYPositionReg_48[9]}},spriteYPositionReg_48}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_48 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1847); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_48 = inSpriteYValue_48[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_48 = $signed(inSpriteYPreScaled_48) >= 11'sh0 & $signed(inSpriteYPreScaled_48) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1450 = {{1{inSpriteYPreScaled_48[10]}},inSpriteYPreScaled_48}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_49 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_49); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_49 = $signed(inSpriteXValue_49) >= 12'sh0 & $signed(inSpriteXValue_49) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1458 = {{1{inSpriteXValue_49[11]}},inSpriteXValue_49}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1849 = {{1{spriteYPositionReg_49[9]}},spriteYPositionReg_49}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_49 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1849); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_49 = inSpriteYValue_49[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_49 = $signed(inSpriteYPreScaled_49) >= 11'sh0 & $signed(inSpriteYPreScaled_49) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1466 = {{1{inSpriteYPreScaled_49[10]}},inSpriteYPreScaled_49}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_50 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_50); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_50 = $signed(inSpriteXValue_50) >= 12'sh0 & $signed(inSpriteXValue_50) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1474 = {{1{inSpriteXValue_50[11]}},inSpriteXValue_50}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1851 = {{1{spriteYPositionReg_50[9]}},spriteYPositionReg_50}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_50 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1851); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_50 = inSpriteYValue_50[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_50 = $signed(inSpriteYPreScaled_50) >= 11'sh0 & $signed(inSpriteYPreScaled_50) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1482 = {{1{inSpriteYPreScaled_50[10]}},inSpriteYPreScaled_50}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_51 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_51); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_51 = $signed(inSpriteXValue_51) >= 12'sh0 & $signed(inSpriteXValue_51) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1490 = {{1{inSpriteXValue_51[11]}},inSpriteXValue_51}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1853 = {{1{spriteYPositionReg_51[9]}},spriteYPositionReg_51}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_51 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1853); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_51 = inSpriteYValue_51[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_51 = $signed(inSpriteYPreScaled_51) >= 11'sh0 & $signed(inSpriteYPreScaled_51) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1498 = {{1{inSpriteYPreScaled_51[10]}},inSpriteYPreScaled_51}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_52 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_52); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_52 = $signed(inSpriteXValue_52) >= 12'sh0 & $signed(inSpriteXValue_52) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1506 = {{1{inSpriteXValue_52[11]}},inSpriteXValue_52}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1855 = {{1{spriteYPositionReg_52[9]}},spriteYPositionReg_52}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_52 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1855); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_52 = inSpriteYValue_52[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_52 = $signed(inSpriteYPreScaled_52) >= 11'sh0 & $signed(inSpriteYPreScaled_52) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1514 = {{1{inSpriteYPreScaled_52[10]}},inSpriteYPreScaled_52}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_53 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_53); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_53 = $signed(inSpriteXValue_53) >= 12'sh0 & $signed(inSpriteXValue_53) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1522 = {{1{inSpriteXValue_53[11]}},inSpriteXValue_53}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1857 = {{1{spriteYPositionReg_53[9]}},spriteYPositionReg_53}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_53 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1857); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_53 = inSpriteYValue_53[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_53 = $signed(inSpriteYPreScaled_53) >= 11'sh0 & $signed(inSpriteYPreScaled_53) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1530 = {{1{inSpriteYPreScaled_53[10]}},inSpriteYPreScaled_53}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_54 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_54); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_54 = $signed(inSpriteXValue_54) >= 12'sh0 & $signed(inSpriteXValue_54) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1538 = {{1{inSpriteXValue_54[11]}},inSpriteXValue_54}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1859 = {{1{spriteYPositionReg_54[9]}},spriteYPositionReg_54}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_54 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1859); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_54 = inSpriteYValue_54[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_54 = $signed(inSpriteYPreScaled_54) >= 11'sh0 & $signed(inSpriteYPreScaled_54) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1546 = {{1{inSpriteYPreScaled_54[10]}},inSpriteYPreScaled_54}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_55 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_55); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_55 = $signed(inSpriteXValue_55) >= 12'sh0 & $signed(inSpriteXValue_55) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1554 = {{1{inSpriteXValue_55[11]}},inSpriteXValue_55}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1861 = {{1{spriteYPositionReg_55[9]}},spriteYPositionReg_55}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_55 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1861); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_55 = inSpriteYValue_55[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_55 = $signed(inSpriteYPreScaled_55) >= 11'sh0 & $signed(inSpriteYPreScaled_55) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1562 = {{1{inSpriteYPreScaled_55[10]}},inSpriteYPreScaled_55}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_56 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_56); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_56 = $signed(inSpriteXValue_56) >= 12'sh0 & $signed(inSpriteXValue_56) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1570 = {{1{inSpriteXValue_56[11]}},inSpriteXValue_56}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1863 = {{1{spriteYPositionReg_56[9]}},spriteYPositionReg_56}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_56 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1863); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_56 = inSpriteYValue_56[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_56 = $signed(inSpriteYPreScaled_56) >= 11'sh0 & $signed(inSpriteYPreScaled_56) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1578 = {{1{inSpriteYPreScaled_56[10]}},inSpriteYPreScaled_56}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_57 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_57); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_57 = $signed(inSpriteXValue_57) >= 12'sh0 & $signed(inSpriteXValue_57) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1586 = {{1{inSpriteXValue_57[11]}},inSpriteXValue_57}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1865 = {{1{spriteYPositionReg_57[9]}},spriteYPositionReg_57}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_57 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1865); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_57 = inSpriteYValue_57[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_57 = $signed(inSpriteYPreScaled_57) >= 11'sh0 & $signed(inSpriteYPreScaled_57) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1594 = {{1{inSpriteYPreScaled_57[10]}},inSpriteYPreScaled_57}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_58 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_58); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_58_T = $signed(inSpriteXValue_58) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_58_T_4 = inSpriteXValue_58[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_58_T_8 = _inSpriteHorizontal_58_T & $signed(inSpriteXValue_58) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_58_T_5 = {$signed(inSpriteXValue_58), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_58_T_14 = _inSpriteHorizontal_58_T & $signed(inSpriteXValue_58) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1600 = spriteScaleUpHorizontalReg_58 ? $signed({{2{_inSpriteX_58_T_4[10]}},_inSpriteX_58_T_4}) :
    $signed(_inSpriteX_58_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1601 = spriteScaleUpHorizontalReg_58 ? _inSpriteHorizontal_58_T_8 : _inSpriteHorizontal_58_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1602 = ~spriteScaleUpHorizontalReg_58 ? $signed({{1{inSpriteXValue_58[11]}},inSpriteXValue_58}) :
    $signed(_GEN_1600); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_58 = ~spriteScaleUpHorizontalReg_58 ? $signed(inSpriteXValue_58) >= 12'sh0 & $signed(
    inSpriteXValue_58) < 12'sh20 : _GEN_1601; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1867 = {{1{spriteYPositionReg_58[9]}},spriteYPositionReg_58}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_58 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1867); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_58 = inSpriteYValue_58[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_58_T = $signed(inSpriteYPreScaled_58) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_58_T_4 = inSpriteYPreScaled_58[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_58_T_8 = _inSpriteVertical_58_T & $signed(inSpriteYPreScaled_58) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_58_T_5 = {$signed(inSpriteYPreScaled_58), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_58_T_14 = _inSpriteVertical_58_T & $signed(inSpriteYPreScaled_58) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1608 = spriteScaleUpVerticalReg_58 ? $signed({{2{_inSpriteY_58_T_4[9]}},_inSpriteY_58_T_4}) :
    $signed(_inSpriteY_58_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1609 = spriteScaleUpVerticalReg_58 ? _inSpriteVertical_58_T_8 : _inSpriteVertical_58_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1610 = ~spriteScaleUpVerticalReg_58 ? $signed({{1{inSpriteYPreScaled_58[10]}},inSpriteYPreScaled_58})
     : $signed(_GEN_1608); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_58 = ~spriteScaleUpVerticalReg_58 ? $signed(inSpriteYPreScaled_58) >= 11'sh0 & $signed(
    inSpriteYPreScaled_58) < 11'sh20 : _GEN_1609; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_59 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_59); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_59_T = $signed(inSpriteXValue_59) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_59_T_4 = inSpriteXValue_59[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_59_T_8 = _inSpriteHorizontal_59_T & $signed(inSpriteXValue_59) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_59_T_5 = {$signed(inSpriteXValue_59), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_59_T_14 = _inSpriteHorizontal_59_T & $signed(inSpriteXValue_59) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1616 = spriteScaleUpHorizontalReg_59 ? $signed({{2{_inSpriteX_59_T_4[10]}},_inSpriteX_59_T_4}) :
    $signed(_inSpriteX_59_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1617 = spriteScaleUpHorizontalReg_59 ? _inSpriteHorizontal_59_T_8 : _inSpriteHorizontal_59_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1618 = ~spriteScaleUpHorizontalReg_59 ? $signed({{1{inSpriteXValue_59[11]}},inSpriteXValue_59}) :
    $signed(_GEN_1616); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_59 = ~spriteScaleUpHorizontalReg_59 ? $signed(inSpriteXValue_59) >= 12'sh0 & $signed(
    inSpriteXValue_59) < 12'sh20 : _GEN_1617; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1869 = {{1{spriteYPositionReg_59[9]}},spriteYPositionReg_59}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_59 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1869); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_59 = inSpriteYValue_59[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_59_T = $signed(inSpriteYPreScaled_59) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_59_T_4 = inSpriteYPreScaled_59[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_59_T_8 = _inSpriteVertical_59_T & $signed(inSpriteYPreScaled_59) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_59_T_5 = {$signed(inSpriteYPreScaled_59), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_59_T_14 = _inSpriteVertical_59_T & $signed(inSpriteYPreScaled_59) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1624 = spriteScaleUpVerticalReg_59 ? $signed({{2{_inSpriteY_59_T_4[9]}},_inSpriteY_59_T_4}) :
    $signed(_inSpriteY_59_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1625 = spriteScaleUpVerticalReg_59 ? _inSpriteVertical_59_T_8 : _inSpriteVertical_59_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1626 = ~spriteScaleUpVerticalReg_59 ? $signed({{1{inSpriteYPreScaled_59[10]}},inSpriteYPreScaled_59})
     : $signed(_GEN_1624); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_59 = ~spriteScaleUpVerticalReg_59 ? $signed(inSpriteYPreScaled_59) >= 11'sh0 & $signed(
    inSpriteYPreScaled_59) < 11'sh20 : _GEN_1625; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_60 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_60); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  _inSpriteHorizontal_60_T = $signed(inSpriteXValue_60) >= 12'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:54]
  wire [10:0] _inSpriteX_60_T_4 = inSpriteXValue_60[11:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 279:47]
  wire  _inSpriteHorizontal_60_T_8 = _inSpriteHorizontal_60_T & $signed(inSpriteXValue_60) < 12'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 280:63]
  wire [12:0] _inSpriteX_60_T_5 = {$signed(inSpriteXValue_60), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 284:45]
  wire  _inSpriteHorizontal_60_T_14 = _inSpriteHorizontal_60_T & $signed(inSpriteXValue_60) < 12'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 288:63]
  wire [12:0] _GEN_1632 = spriteScaleUpHorizontalReg_60 ? $signed({{2{_inSpriteX_60_T_4[10]}},_inSpriteX_60_T_4}) :
    $signed(_inSpriteX_60_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48 284:20]
  wire  _GEN_1633 = spriteScaleUpHorizontalReg_60 ? _inSpriteHorizontal_60_T_8 : _inSpriteHorizontal_60_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 273:48]
  wire [12:0] _GEN_1634 = ~spriteScaleUpHorizontalReg_60 ? $signed({{1{inSpriteXValue_60[11]}},inSpriteXValue_60}) :
    $signed(_GEN_1632); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire  inSpriteHorizontal_60 = ~spriteScaleUpHorizontalReg_60 ? $signed(inSpriteXValue_60) >= 12'sh0 & $signed(
    inSpriteXValue_60) < 12'sh20 : _GEN_1633; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 272:29]
  wire [10:0] _GEN_1871 = {{1{spriteYPositionReg_60[9]}},spriteYPositionReg_60}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_60 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1871); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_60 = inSpriteYValue_60[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  _inSpriteVertical_60_T = $signed(inSpriteYPreScaled_60) >= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:52]
  wire [9:0] _inSpriteY_60_T_4 = inSpriteYPreScaled_60[10:1]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 308:47]
  wire  _inSpriteVertical_60_T_8 = _inSpriteVertical_60_T & $signed(inSpriteYPreScaled_60) < 11'sh40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 309:61]
  wire [11:0] _inSpriteY_60_T_5 = {$signed(inSpriteYPreScaled_60), 1'h0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 313:45]
  wire  _inSpriteVertical_60_T_14 = _inSpriteVertical_60_T & $signed(inSpriteYPreScaled_60) < 11'sh10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 317:61]
  wire [11:0] _GEN_1640 = spriteScaleUpVerticalReg_60 ? $signed({{2{_inSpriteY_60_T_4[9]}},_inSpriteY_60_T_4}) :
    $signed(_inSpriteY_60_T_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45 313:20]
  wire  _GEN_1641 = spriteScaleUpVerticalReg_60 ? _inSpriteVertical_60_T_8 : _inSpriteVertical_60_T_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 302:45]
  wire [11:0] _GEN_1642 = ~spriteScaleUpVerticalReg_60 ? $signed({{1{inSpriteYPreScaled_60[10]}},inSpriteYPreScaled_60})
     : $signed(_GEN_1640); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire  inSpriteVertical_60 = ~spriteScaleUpVerticalReg_60 ? $signed(inSpriteYPreScaled_60) >= 11'sh0 & $signed(
    inSpriteYPreScaled_60) < 11'sh20 : _GEN_1641; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 301:27]
  wire [11:0] inSpriteXValue_61 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_61); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_61 = $signed(inSpriteXValue_61) >= 12'sh0 & $signed(inSpriteXValue_61) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1650 = {{1{inSpriteXValue_61[11]}},inSpriteXValue_61}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1873 = {{1{spriteYPositionReg_61[9]}},spriteYPositionReg_61}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_61 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1873); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_61 = inSpriteYValue_61[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_61 = $signed(inSpriteYPreScaled_61) >= 11'sh0 & $signed(inSpriteYPreScaled_61) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1658 = {{1{inSpriteYPreScaled_61[10]}},inSpriteYPreScaled_61}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_62 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_62); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_62 = $signed(inSpriteXValue_62) >= 12'sh0 & $signed(inSpriteXValue_62) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1666 = {{1{inSpriteXValue_62[11]}},inSpriteXValue_62}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1875 = {{1{spriteYPositionReg_62[9]}},spriteYPositionReg_62}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_62 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1875); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_62 = inSpriteYValue_62[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_62 = $signed(inSpriteYPreScaled_62) >= 11'sh0 & $signed(inSpriteYPreScaled_62) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1674 = {{1{inSpriteYPreScaled_62[10]}},inSpriteYPreScaled_62}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_63 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_63); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_63 = $signed(inSpriteXValue_63) >= 12'sh0 & $signed(inSpriteXValue_63) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_1682 = {{1{inSpriteXValue_63[11]}},inSpriteXValue_63}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_1877 = {{1{spriteYPositionReg_63[9]}},spriteYPositionReg_63}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_63 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_1877); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_63 = inSpriteYValue_63[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_63 = $signed(inSpriteYPreScaled_63) >= 11'sh0 & $signed(inSpriteYPreScaled_63) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_1690 = {{1{inSpriteYPreScaled_63[10]}},inSpriteYPreScaled_63}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteX_0 = _GEN_674[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_0 = _GEN_682[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_0_io_address_T_2 = 6'h20 * inSpriteY_0[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1881 = {{6'd0}, inSpriteX_0[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_0_io_address_T_4 = _GEN_1881 + _spriteMemories_0_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_3 = _GEN_722[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_3 = _GEN_730[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_3_io_address_T_2 = 6'h20 * inSpriteY_3[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1890 = {{6'd0}, inSpriteX_3[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_3_io_address_T_4 = _GEN_1890 + _spriteMemories_3_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_7 = _GEN_786[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_7 = _GEN_794[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_7_io_address_T_2 = 6'h20 * inSpriteY_7[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1902 = {{6'd0}, inSpriteX_7[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_7_io_address_T_4 = _GEN_1902 + _spriteMemories_7_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_8 = _GEN_802[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_8 = _GEN_810[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_8_io_address_T_2 = 6'h20 * inSpriteY_8[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1905 = {{6'd0}, inSpriteX_8[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_8_io_address_T_4 = _GEN_1905 + _spriteMemories_8_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_9 = _GEN_818[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_9 = _GEN_826[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_9_io_address_T_2 = 6'h20 * inSpriteY_9[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1908 = {{6'd0}, inSpriteX_9[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_9_io_address_T_4 = _GEN_1908 + _spriteMemories_9_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_10 = _GEN_834[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_10 = _GEN_842[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_10_io_address_T_2 = 6'h20 * inSpriteY_10[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1911 = {{6'd0}, inSpriteX_10[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_10_io_address_T_4 = _GEN_1911 + _spriteMemories_10_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_11 = _GEN_850[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_11 = _GEN_858[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_11_io_address_T_2 = 6'h20 * inSpriteY_11[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1914 = {{6'd0}, inSpriteX_11[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_11_io_address_T_4 = _GEN_1914 + _spriteMemories_11_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_12 = _GEN_866[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_12 = _GEN_874[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_12_io_address_T_2 = 6'h20 * inSpriteY_12[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1917 = {{6'd0}, inSpriteX_12[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_12_io_address_T_4 = _GEN_1917 + _spriteMemories_12_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_13 = _GEN_882[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_13 = _GEN_890[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_13_io_address_T_2 = 6'h20 * inSpriteY_13[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1920 = {{6'd0}, inSpriteX_13[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_13_io_address_T_4 = _GEN_1920 + _spriteMemories_13_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_14 = _GEN_898[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_14 = _GEN_906[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_14_io_address_T_2 = 6'h20 * inSpriteY_14[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1923 = {{6'd0}, inSpriteX_14[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_14_io_address_T_4 = _GEN_1923 + _spriteMemories_14_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_16 = _GEN_930[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_16 = _GEN_938[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_16_io_address_T_2 = 6'h20 * inSpriteY_16[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1929 = {{6'd0}, inSpriteX_16[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_16_io_address_T_4 = _GEN_1929 + _spriteMemories_16_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_17 = _GEN_946[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_17 = _GEN_954[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_17_io_address_T_2 = 6'h20 * inSpriteY_17[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1932 = {{6'd0}, inSpriteX_17[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_17_io_address_T_4 = _GEN_1932 + _spriteMemories_17_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_18 = _GEN_962[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_18 = _GEN_970[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_18_io_address_T_2 = 6'h20 * inSpriteY_18[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1935 = {{6'd0}, inSpriteX_18[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_18_io_address_T_4 = _GEN_1935 + _spriteMemories_18_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_19 = _GEN_978[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_19 = _GEN_986[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_19_io_address_T_2 = 6'h20 * inSpriteY_19[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1938 = {{6'd0}, inSpriteX_19[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_19_io_address_T_4 = _GEN_1938 + _spriteMemories_19_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_20 = _GEN_994[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_20 = _GEN_1002[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_20_io_address_T_2 = 6'h20 * inSpriteY_20[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1941 = {{6'd0}, inSpriteX_20[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_20_io_address_T_4 = _GEN_1941 + _spriteMemories_20_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_21 = _GEN_1010[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_21 = _GEN_1018[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_21_io_address_T_2 = 6'h20 * inSpriteY_21[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1944 = {{6'd0}, inSpriteX_21[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_21_io_address_T_4 = _GEN_1944 + _spriteMemories_21_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_22 = _GEN_1026[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_22 = _GEN_1034[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_22_io_address_T_2 = 6'h20 * inSpriteY_22[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1947 = {{6'd0}, inSpriteX_22[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_22_io_address_T_4 = _GEN_1947 + _spriteMemories_22_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_23 = _GEN_1042[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_23 = _GEN_1050[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_23_io_address_T_2 = 6'h20 * inSpriteY_23[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1950 = {{6'd0}, inSpriteX_23[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_23_io_address_T_4 = _GEN_1950 + _spriteMemories_23_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_24 = _GEN_1058[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_24 = _GEN_1066[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_24_io_address_T_2 = 6'h20 * inSpriteY_24[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1953 = {{6'd0}, inSpriteX_24[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_24_io_address_T_4 = _GEN_1953 + _spriteMemories_24_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_25 = _GEN_1074[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_25 = _GEN_1082[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_25_io_address_T_2 = 6'h20 * inSpriteY_25[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1956 = {{6'd0}, inSpriteX_25[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_25_io_address_T_4 = _GEN_1956 + _spriteMemories_25_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_26 = _GEN_1090[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_26 = _GEN_1098[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_26_io_address_T_2 = 6'h20 * inSpriteY_26[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1959 = {{6'd0}, inSpriteX_26[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_26_io_address_T_4 = _GEN_1959 + _spriteMemories_26_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_27 = _GEN_1106[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_27 = _GEN_1114[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_27_io_address_T_2 = 6'h20 * inSpriteY_27[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1962 = {{6'd0}, inSpriteX_27[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_27_io_address_T_4 = _GEN_1962 + _spriteMemories_27_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_28 = _GEN_1122[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_28 = _GEN_1130[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_28_io_address_T_2 = 6'h20 * inSpriteY_28[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1965 = {{6'd0}, inSpriteX_28[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_28_io_address_T_4 = _GEN_1965 + _spriteMemories_28_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_29 = _GEN_1138[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_29 = _GEN_1146[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_29_io_address_T_2 = 6'h20 * inSpriteY_29[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1968 = {{6'd0}, inSpriteX_29[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_29_io_address_T_4 = _GEN_1968 + _spriteMemories_29_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_30 = _GEN_1154[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_30 = _GEN_1162[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_30_io_address_T_2 = 6'h20 * inSpriteY_30[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1971 = {{6'd0}, inSpriteX_30[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_30_io_address_T_4 = _GEN_1971 + _spriteMemories_30_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_31 = _GEN_1170[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_31 = _GEN_1178[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_31_io_address_T_2 = 6'h20 * inSpriteY_31[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1974 = {{6'd0}, inSpriteX_31[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_31_io_address_T_4 = _GEN_1974 + _spriteMemories_31_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_32 = _GEN_1186[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_32 = _GEN_1194[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_32_io_address_T_2 = 6'h20 * inSpriteY_32[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1977 = {{6'd0}, inSpriteX_32[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_32_io_address_T_4 = _GEN_1977 + _spriteMemories_32_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_33 = _GEN_1202[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_33 = _GEN_1210[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_33_io_address_T_2 = 6'h20 * inSpriteY_33[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1980 = {{6'd0}, inSpriteX_33[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_33_io_address_T_4 = _GEN_1980 + _spriteMemories_33_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_34 = _GEN_1218[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_34 = _GEN_1226[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_34_io_address_T_2 = 6'h20 * inSpriteY_34[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1983 = {{6'd0}, inSpriteX_34[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_34_io_address_T_4 = _GEN_1983 + _spriteMemories_34_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_35 = _GEN_1234[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_35 = _GEN_1242[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_35_io_address_T_2 = 6'h20 * inSpriteY_35[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1986 = {{6'd0}, inSpriteX_35[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_35_io_address_T_4 = _GEN_1986 + _spriteMemories_35_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_36 = _GEN_1250[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_36 = _GEN_1258[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_36_io_address_T_2 = 6'h20 * inSpriteY_36[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1989 = {{6'd0}, inSpriteX_36[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_36_io_address_T_4 = _GEN_1989 + _spriteMemories_36_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_37 = _GEN_1266[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_37 = _GEN_1274[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_37_io_address_T_2 = 6'h20 * inSpriteY_37[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1992 = {{6'd0}, inSpriteX_37[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_37_io_address_T_4 = _GEN_1992 + _spriteMemories_37_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_38 = _GEN_1282[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_38 = _GEN_1290[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_38_io_address_T_2 = 6'h20 * inSpriteY_38[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1995 = {{6'd0}, inSpriteX_38[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_38_io_address_T_4 = _GEN_1995 + _spriteMemories_38_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_39 = _GEN_1298[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_39 = _GEN_1306[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_39_io_address_T_2 = 6'h20 * inSpriteY_39[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1998 = {{6'd0}, inSpriteX_39[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_39_io_address_T_4 = _GEN_1998 + _spriteMemories_39_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_40 = _GEN_1314[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_40 = _GEN_1322[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_40_io_address_T_2 = 6'h20 * inSpriteY_40[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2001 = {{6'd0}, inSpriteX_40[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_40_io_address_T_4 = _GEN_2001 + _spriteMemories_40_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_41 = _GEN_1330[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_41 = _GEN_1338[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_41_io_address_T_2 = 6'h20 * inSpriteY_41[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2004 = {{6'd0}, inSpriteX_41[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_41_io_address_T_4 = _GEN_2004 + _spriteMemories_41_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_42 = _GEN_1346[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_42 = _GEN_1354[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_42_io_address_T_2 = 6'h20 * inSpriteY_42[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2007 = {{6'd0}, inSpriteX_42[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_42_io_address_T_4 = _GEN_2007 + _spriteMemories_42_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_43 = _GEN_1362[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_43 = _GEN_1370[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_43_io_address_T_2 = 6'h20 * inSpriteY_43[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2010 = {{6'd0}, inSpriteX_43[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_43_io_address_T_4 = _GEN_2010 + _spriteMemories_43_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_44 = _GEN_1378[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_44 = _GEN_1386[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_44_io_address_T_2 = 6'h20 * inSpriteY_44[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2013 = {{6'd0}, inSpriteX_44[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_44_io_address_T_4 = _GEN_2013 + _spriteMemories_44_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_45 = _GEN_1394[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_45 = _GEN_1402[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_45_io_address_T_2 = 6'h20 * inSpriteY_45[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2016 = {{6'd0}, inSpriteX_45[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_45_io_address_T_4 = _GEN_2016 + _spriteMemories_45_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_46 = _GEN_1410[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_46 = _GEN_1418[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_46_io_address_T_2 = 6'h20 * inSpriteY_46[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2019 = {{6'd0}, inSpriteX_46[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_46_io_address_T_4 = _GEN_2019 + _spriteMemories_46_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_47 = _GEN_1426[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_47 = _GEN_1434[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_47_io_address_T_2 = 6'h20 * inSpriteY_47[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2022 = {{6'd0}, inSpriteX_47[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_47_io_address_T_4 = _GEN_2022 + _spriteMemories_47_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_48 = _GEN_1442[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_48 = _GEN_1450[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_48_io_address_T_2 = 6'h20 * inSpriteY_48[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2025 = {{6'd0}, inSpriteX_48[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_48_io_address_T_4 = _GEN_2025 + _spriteMemories_48_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_49 = _GEN_1458[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_49 = _GEN_1466[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_49_io_address_T_2 = 6'h20 * inSpriteY_49[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2028 = {{6'd0}, inSpriteX_49[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_49_io_address_T_4 = _GEN_2028 + _spriteMemories_49_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_50 = _GEN_1474[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_50 = _GEN_1482[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_50_io_address_T_2 = 6'h20 * inSpriteY_50[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2031 = {{6'd0}, inSpriteX_50[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_50_io_address_T_4 = _GEN_2031 + _spriteMemories_50_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_51 = _GEN_1490[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_51 = _GEN_1498[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_51_io_address_T_2 = 6'h20 * inSpriteY_51[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2034 = {{6'd0}, inSpriteX_51[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_51_io_address_T_4 = _GEN_2034 + _spriteMemories_51_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_52 = _GEN_1506[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_52 = _GEN_1514[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_52_io_address_T_2 = 6'h20 * inSpriteY_52[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2037 = {{6'd0}, inSpriteX_52[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_52_io_address_T_4 = _GEN_2037 + _spriteMemories_52_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_53 = _GEN_1522[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_53 = _GEN_1530[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_53_io_address_T_2 = 6'h20 * inSpriteY_53[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2040 = {{6'd0}, inSpriteX_53[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_53_io_address_T_4 = _GEN_2040 + _spriteMemories_53_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_54 = _GEN_1538[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_54 = _GEN_1546[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_54_io_address_T_2 = 6'h20 * inSpriteY_54[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2043 = {{6'd0}, inSpriteX_54[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_54_io_address_T_4 = _GEN_2043 + _spriteMemories_54_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_55 = _GEN_1554[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_55 = _GEN_1562[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_55_io_address_T_2 = 6'h20 * inSpriteY_55[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2046 = {{6'd0}, inSpriteX_55[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_55_io_address_T_4 = _GEN_2046 + _spriteMemories_55_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_56 = _GEN_1570[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_56 = _GEN_1578[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_56_io_address_T_2 = 6'h20 * inSpriteY_56[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2049 = {{6'd0}, inSpriteX_56[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_56_io_address_T_4 = _GEN_2049 + _spriteMemories_56_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_57 = _GEN_1586[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_57 = _GEN_1594[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_57_io_address_T_2 = 6'h20 * inSpriteY_57[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2052 = {{6'd0}, inSpriteX_57[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_57_io_address_T_4 = _GEN_2052 + _spriteMemories_57_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_58 = _GEN_1602[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_58 = _GEN_1610[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_58_io_address_T_2 = 6'h20 * inSpriteY_58[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2055 = {{6'd0}, inSpriteX_58[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_58_io_address_T_4 = _GEN_2055 + _spriteMemories_58_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_59 = _GEN_1618[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_59 = _GEN_1626[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_59_io_address_T_2 = 6'h20 * inSpriteY_59[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2058 = {{6'd0}, inSpriteX_59[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_59_io_address_T_4 = _GEN_2058 + _spriteMemories_59_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_60 = _GEN_1634[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_60 = _GEN_1642[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_60_io_address_T_2 = 6'h20 * inSpriteY_60[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2061 = {{6'd0}, inSpriteX_60[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_60_io_address_T_4 = _GEN_2061 + _spriteMemories_60_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_61 = _GEN_1650[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_61 = _GEN_1658[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_61_io_address_T_2 = 6'h20 * inSpriteY_61[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2064 = {{6'd0}, inSpriteX_61[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_61_io_address_T_4 = _GEN_2064 + _spriteMemories_61_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_62 = _GEN_1666[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_62 = _GEN_1674[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_62_io_address_T_2 = 6'h20 * inSpriteY_62[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2067 = {{6'd0}, inSpriteX_62[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_62_io_address_T_4 = _GEN_2067 + _spriteMemories_62_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_63 = _GEN_1682[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_63 = _GEN_1690[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_63_io_address_T_2 = 6'h20 * inSpriteY_63[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_2070 = {{6'd0}, inSpriteX_63[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_63_io_address_T_4 = _GEN_2070 + _spriteMemories_63_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] pixelColorSprite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 339:33]
  reg  pixelColorSpriteValid; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 340:38]
  wire [5:0] pixelColorInDisplay = pixelColorSpriteValid ? pixelColorSprite : pixelColorBack; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 344:32]
  reg  pixelColourVGA_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  pixelColourVGA_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  pixelColourVGA_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  wire [5:0] pixelColourVGA = pixelColourVGA_pipeReg_0 ? pixelColorInDisplay : 6'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 345:27]
  reg [3:0] io_vgaRed_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 349:23]
  reg [3:0] io_vgaGreen_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 350:25]
  reg [3:0] io_vgaBlue_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 351:24]
  Memory backTileMemories_0 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_0_clock),
    .io_address(backTileMemories_0_io_address),
    .io_dataRead(backTileMemories_0_io_dataRead)
  );
  Memory_1 backTileMemories_1 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_1_clock),
    .io_address(backTileMemories_1_io_address),
    .io_dataRead(backTileMemories_1_io_dataRead)
  );
  Memory_2 backTileMemories_2 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_2_clock),
    .io_address(backTileMemories_2_io_address),
    .io_dataRead(backTileMemories_2_io_dataRead)
  );
  Memory_3 backTileMemories_3 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_3_clock),
    .io_address(backTileMemories_3_io_address),
    .io_dataRead(backTileMemories_3_io_dataRead)
  );
  Memory_4 backTileMemories_4 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_4_clock),
    .io_address(backTileMemories_4_io_address),
    .io_dataRead(backTileMemories_4_io_dataRead)
  );
  Memory_5 backTileMemories_5 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_5_clock),
    .io_address(backTileMemories_5_io_address),
    .io_dataRead(backTileMemories_5_io_dataRead)
  );
  Memory_6 backTileMemories_6 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_6_clock),
    .io_address(backTileMemories_6_io_address),
    .io_dataRead(backTileMemories_6_io_dataRead)
  );
  Memory_7 backTileMemories_7 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_7_clock),
    .io_address(backTileMemories_7_io_address),
    .io_dataRead(backTileMemories_7_io_dataRead)
  );
  Memory_8 backTileMemories_8 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_8_clock),
    .io_address(backTileMemories_8_io_address),
    .io_dataRead(backTileMemories_8_io_dataRead)
  );
  Memory_9 backTileMemories_9 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_9_clock),
    .io_address(backTileMemories_9_io_address),
    .io_dataRead(backTileMemories_9_io_dataRead)
  );
  Memory_10 backTileMemories_10 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_10_clock),
    .io_address(backTileMemories_10_io_address),
    .io_dataRead(backTileMemories_10_io_dataRead)
  );
  Memory_11 backTileMemories_11 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_11_clock),
    .io_address(backTileMemories_11_io_address),
    .io_dataRead(backTileMemories_11_io_dataRead)
  );
  Memory_12 backTileMemories_12 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_12_clock),
    .io_address(backTileMemories_12_io_address),
    .io_dataRead(backTileMemories_12_io_dataRead)
  );
  Memory_13 backTileMemories_13 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_13_clock),
    .io_address(backTileMemories_13_io_address),
    .io_dataRead(backTileMemories_13_io_dataRead)
  );
  Memory_14 backTileMemories_14 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_14_clock),
    .io_address(backTileMemories_14_io_address),
    .io_dataRead(backTileMemories_14_io_dataRead)
  );
  Memory_15 backTileMemories_15 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_15_clock),
    .io_address(backTileMemories_15_io_address),
    .io_dataRead(backTileMemories_15_io_dataRead)
  );
  Memory_16 backTileMemories_16 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_16_clock),
    .io_address(backTileMemories_16_io_address),
    .io_dataRead(backTileMemories_16_io_dataRead)
  );
  Memory_17 backTileMemories_17 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_17_clock),
    .io_address(backTileMemories_17_io_address),
    .io_dataRead(backTileMemories_17_io_dataRead)
  );
  Memory_18 backTileMemories_18 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_18_clock),
    .io_address(backTileMemories_18_io_address),
    .io_dataRead(backTileMemories_18_io_dataRead)
  );
  Memory_19 backTileMemories_19 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_19_clock),
    .io_address(backTileMemories_19_io_address),
    .io_dataRead(backTileMemories_19_io_dataRead)
  );
  Memory_20 backTileMemories_20 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_20_clock),
    .io_address(backTileMemories_20_io_address),
    .io_dataRead(backTileMemories_20_io_dataRead)
  );
  Memory_21 backTileMemories_21 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_21_clock),
    .io_address(backTileMemories_21_io_address),
    .io_dataRead(backTileMemories_21_io_dataRead)
  );
  Memory_22 backTileMemories_22 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_22_clock),
    .io_address(backTileMemories_22_io_address),
    .io_dataRead(backTileMemories_22_io_dataRead)
  );
  Memory_23 backTileMemories_23 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_23_clock),
    .io_address(backTileMemories_23_io_address),
    .io_dataRead(backTileMemories_23_io_dataRead)
  );
  Memory_24 backTileMemories_24 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_24_clock),
    .io_address(backTileMemories_24_io_address),
    .io_dataRead(backTileMemories_24_io_dataRead)
  );
  Memory_25 backTileMemories_25 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_25_clock),
    .io_address(backTileMemories_25_io_address),
    .io_dataRead(backTileMemories_25_io_dataRead)
  );
  Memory_26 backTileMemories_26 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_26_clock),
    .io_address(backTileMemories_26_io_address),
    .io_dataRead(backTileMemories_26_io_dataRead)
  );
  Memory_27 backTileMemories_27 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_27_clock),
    .io_address(backTileMemories_27_io_address),
    .io_dataRead(backTileMemories_27_io_dataRead)
  );
  Memory_28 backTileMemories_28 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_28_clock),
    .io_address(backTileMemories_28_io_address),
    .io_dataRead(backTileMemories_28_io_dataRead)
  );
  Memory_29 backTileMemories_29 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_29_clock),
    .io_address(backTileMemories_29_io_address),
    .io_dataRead(backTileMemories_29_io_dataRead)
  );
  Memory_30 backTileMemories_30 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_30_clock),
    .io_address(backTileMemories_30_io_address),
    .io_dataRead(backTileMemories_30_io_dataRead)
  );
  Memory_31 backTileMemories_31 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_31_clock),
    .io_address(backTileMemories_31_io_address),
    .io_dataRead(backTileMemories_31_io_dataRead)
  );
  Memory_32 backTileMemories_32 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_32_clock),
    .io_address(backTileMemories_32_io_address),
    .io_dataRead(backTileMemories_32_io_dataRead)
  );
  Memory_33 backTileMemories_33 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_33_clock),
    .io_address(backTileMemories_33_io_address),
    .io_dataRead(backTileMemories_33_io_dataRead)
  );
  Memory_34 backTileMemories_34 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_34_clock),
    .io_address(backTileMemories_34_io_address),
    .io_dataRead(backTileMemories_34_io_dataRead)
  );
  Memory_35 backTileMemories_35 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_35_clock),
    .io_address(backTileMemories_35_io_address),
    .io_dataRead(backTileMemories_35_io_dataRead)
  );
  Memory_36 backTileMemories_36 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_36_clock),
    .io_address(backTileMemories_36_io_address),
    .io_dataRead(backTileMemories_36_io_dataRead)
  );
  Memory_37 backTileMemories_37 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_37_clock),
    .io_address(backTileMemories_37_io_address),
    .io_dataRead(backTileMemories_37_io_dataRead)
  );
  Memory_38 backTileMemories_38 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_38_clock),
    .io_address(backTileMemories_38_io_address),
    .io_dataRead(backTileMemories_38_io_dataRead)
  );
  Memory_39 backTileMemories_39 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_39_clock),
    .io_address(backTileMemories_39_io_address),
    .io_dataRead(backTileMemories_39_io_dataRead)
  );
  Memory_40 backTileMemories_40 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_40_clock),
    .io_address(backTileMemories_40_io_address),
    .io_dataRead(backTileMemories_40_io_dataRead)
  );
  Memory_41 backTileMemories_41 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_41_clock),
    .io_address(backTileMemories_41_io_address),
    .io_dataRead(backTileMemories_41_io_dataRead)
  );
  Memory_42 backTileMemories_42 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_42_clock),
    .io_address(backTileMemories_42_io_address),
    .io_dataRead(backTileMemories_42_io_dataRead)
  );
  Memory_43 backTileMemories_43 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_43_clock),
    .io_address(backTileMemories_43_io_address),
    .io_dataRead(backTileMemories_43_io_dataRead)
  );
  Memory_44 backTileMemories_44 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_44_clock),
    .io_address(backTileMemories_44_io_address),
    .io_dataRead(backTileMemories_44_io_dataRead)
  );
  Memory_45 backTileMemories_45 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_45_clock),
    .io_address(backTileMemories_45_io_address),
    .io_dataRead(backTileMemories_45_io_dataRead)
  );
  Memory_46 backTileMemories_46 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_46_clock),
    .io_address(backTileMemories_46_io_address),
    .io_dataRead(backTileMemories_46_io_dataRead)
  );
  Memory_47 backTileMemories_47 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_47_clock),
    .io_address(backTileMemories_47_io_address),
    .io_dataRead(backTileMemories_47_io_dataRead)
  );
  Memory_48 backTileMemories_48 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_48_clock),
    .io_address(backTileMemories_48_io_address),
    .io_dataRead(backTileMemories_48_io_dataRead)
  );
  Memory_49 backTileMemories_49 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_49_clock),
    .io_address(backTileMemories_49_io_address),
    .io_dataRead(backTileMemories_49_io_dataRead)
  );
  Memory_50 backTileMemories_50 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_50_clock),
    .io_address(backTileMemories_50_io_address),
    .io_dataRead(backTileMemories_50_io_dataRead)
  );
  Memory_51 backTileMemories_51 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_51_clock),
    .io_address(backTileMemories_51_io_address),
    .io_dataRead(backTileMemories_51_io_dataRead)
  );
  Memory_52 backTileMemories_52 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_52_clock),
    .io_address(backTileMemories_52_io_address),
    .io_dataRead(backTileMemories_52_io_dataRead)
  );
  Memory_53 backTileMemories_53 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_53_clock),
    .io_address(backTileMemories_53_io_address),
    .io_dataRead(backTileMemories_53_io_dataRead)
  );
  Memory_54 backTileMemories_54 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_54_clock),
    .io_address(backTileMemories_54_io_address),
    .io_dataRead(backTileMemories_54_io_dataRead)
  );
  Memory_55 backTileMemories_55 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_55_clock),
    .io_address(backTileMemories_55_io_address),
    .io_dataRead(backTileMemories_55_io_dataRead)
  );
  Memory_56 backTileMemories_56 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_56_clock),
    .io_address(backTileMemories_56_io_address),
    .io_dataRead(backTileMemories_56_io_dataRead)
  );
  Memory_57 backTileMemories_57 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_57_clock),
    .io_address(backTileMemories_57_io_address),
    .io_dataRead(backTileMemories_57_io_dataRead)
  );
  Memory_58 backTileMemories_58 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_58_clock),
    .io_address(backTileMemories_58_io_address),
    .io_dataRead(backTileMemories_58_io_dataRead)
  );
  Memory_59 backTileMemories_59 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_59_clock),
    .io_address(backTileMemories_59_io_address),
    .io_dataRead(backTileMemories_59_io_dataRead)
  );
  Memory_60 backTileMemories_60 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_60_clock),
    .io_address(backTileMemories_60_io_address),
    .io_dataRead(backTileMemories_60_io_dataRead)
  );
  Memory_61 backTileMemories_61 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_61_clock),
    .io_address(backTileMemories_61_io_address),
    .io_dataRead(backTileMemories_61_io_dataRead)
  );
  Memory_62 backTileMemories_62 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_62_clock),
    .io_address(backTileMemories_62_io_address),
    .io_dataRead(backTileMemories_62_io_dataRead)
  );
  Memory_63 backTileMemories_63 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_63_clock),
    .io_address(backTileMemories_63_io_address),
    .io_dataRead(backTileMemories_63_io_dataRead)
  );
  Memory_64 backBufferMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
    .clock(backBufferMemory_clock),
    .io_address(backBufferMemory_io_address),
    .io_dataRead(backBufferMemory_io_dataRead),
    .io_writeEnable(backBufferMemory_io_writeEnable),
    .io_dataWrite(backBufferMemory_io_dataWrite)
  );
  Memory_64 backBufferShadowMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
    .clock(backBufferShadowMemory_clock),
    .io_address(backBufferShadowMemory_io_address),
    .io_dataRead(backBufferShadowMemory_io_dataRead),
    .io_writeEnable(backBufferShadowMemory_io_writeEnable),
    .io_dataWrite(backBufferShadowMemory_io_dataWrite)
  );
  Memory_66 backBufferRestoreMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
    .clock(backBufferRestoreMemory_clock),
    .io_address(backBufferRestoreMemory_io_address),
    .io_dataRead(backBufferRestoreMemory_io_dataRead)
  );
  Memory_67 spriteMemories_0 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_0_clock),
    .io_address(spriteMemories_0_io_address),
    .io_dataRead(spriteMemories_0_io_dataRead)
  );
  Memory_68 spriteMemories_1 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_1_clock),
    .io_address(spriteMemories_1_io_address),
    .io_dataRead(spriteMemories_1_io_dataRead)
  );
  Memory_69 spriteMemories_2 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_2_clock),
    .io_address(spriteMemories_2_io_address),
    .io_dataRead(spriteMemories_2_io_dataRead)
  );
  Memory_70 spriteMemories_3 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_3_clock),
    .io_address(spriteMemories_3_io_address),
    .io_dataRead(spriteMemories_3_io_dataRead)
  );
  Memory_71 spriteMemories_4 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_4_clock),
    .io_address(spriteMemories_4_io_address),
    .io_dataRead(spriteMemories_4_io_dataRead)
  );
  Memory_72 spriteMemories_5 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_5_clock),
    .io_address(spriteMemories_5_io_address),
    .io_dataRead(spriteMemories_5_io_dataRead)
  );
  Memory_73 spriteMemories_6 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_6_clock),
    .io_address(spriteMemories_6_io_address),
    .io_dataRead(spriteMemories_6_io_dataRead)
  );
  Memory_74 spriteMemories_7 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_7_clock),
    .io_address(spriteMemories_7_io_address),
    .io_dataRead(spriteMemories_7_io_dataRead)
  );
  Memory_75 spriteMemories_8 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_8_clock),
    .io_address(spriteMemories_8_io_address),
    .io_dataRead(spriteMemories_8_io_dataRead)
  );
  Memory_76 spriteMemories_9 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_9_clock),
    .io_address(spriteMemories_9_io_address),
    .io_dataRead(spriteMemories_9_io_dataRead)
  );
  Memory_77 spriteMemories_10 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_10_clock),
    .io_address(spriteMemories_10_io_address),
    .io_dataRead(spriteMemories_10_io_dataRead)
  );
  Memory_78 spriteMemories_11 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_11_clock),
    .io_address(spriteMemories_11_io_address),
    .io_dataRead(spriteMemories_11_io_dataRead)
  );
  Memory_79 spriteMemories_12 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_12_clock),
    .io_address(spriteMemories_12_io_address),
    .io_dataRead(spriteMemories_12_io_dataRead)
  );
  Memory_80 spriteMemories_13 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_13_clock),
    .io_address(spriteMemories_13_io_address),
    .io_dataRead(spriteMemories_13_io_dataRead)
  );
  Memory_81 spriteMemories_14 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_14_clock),
    .io_address(spriteMemories_14_io_address),
    .io_dataRead(spriteMemories_14_io_dataRead)
  );
  Memory_82 spriteMemories_15 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_15_clock),
    .io_address(spriteMemories_15_io_address),
    .io_dataRead(spriteMemories_15_io_dataRead)
  );
  Memory_83 spriteMemories_16 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_16_clock),
    .io_address(spriteMemories_16_io_address),
    .io_dataRead(spriteMemories_16_io_dataRead)
  );
  Memory_84 spriteMemories_17 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_17_clock),
    .io_address(spriteMemories_17_io_address),
    .io_dataRead(spriteMemories_17_io_dataRead)
  );
  Memory_85 spriteMemories_18 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_18_clock),
    .io_address(spriteMemories_18_io_address),
    .io_dataRead(spriteMemories_18_io_dataRead)
  );
  Memory_86 spriteMemories_19 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_19_clock),
    .io_address(spriteMemories_19_io_address),
    .io_dataRead(spriteMemories_19_io_dataRead)
  );
  Memory_87 spriteMemories_20 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_20_clock),
    .io_address(spriteMemories_20_io_address),
    .io_dataRead(spriteMemories_20_io_dataRead)
  );
  Memory_88 spriteMemories_21 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_21_clock),
    .io_address(spriteMemories_21_io_address),
    .io_dataRead(spriteMemories_21_io_dataRead)
  );
  Memory_89 spriteMemories_22 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_22_clock),
    .io_address(spriteMemories_22_io_address),
    .io_dataRead(spriteMemories_22_io_dataRead)
  );
  Memory_90 spriteMemories_23 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_23_clock),
    .io_address(spriteMemories_23_io_address),
    .io_dataRead(spriteMemories_23_io_dataRead)
  );
  Memory_91 spriteMemories_24 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_24_clock),
    .io_address(spriteMemories_24_io_address),
    .io_dataRead(spriteMemories_24_io_dataRead)
  );
  Memory_92 spriteMemories_25 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_25_clock),
    .io_address(spriteMemories_25_io_address),
    .io_dataRead(spriteMemories_25_io_dataRead)
  );
  Memory_93 spriteMemories_26 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_26_clock),
    .io_address(spriteMemories_26_io_address),
    .io_dataRead(spriteMemories_26_io_dataRead)
  );
  Memory_94 spriteMemories_27 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_27_clock),
    .io_address(spriteMemories_27_io_address),
    .io_dataRead(spriteMemories_27_io_dataRead)
  );
  Memory_95 spriteMemories_28 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_28_clock),
    .io_address(spriteMemories_28_io_address),
    .io_dataRead(spriteMemories_28_io_dataRead)
  );
  Memory_96 spriteMemories_29 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_29_clock),
    .io_address(spriteMemories_29_io_address),
    .io_dataRead(spriteMemories_29_io_dataRead)
  );
  Memory_97 spriteMemories_30 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_30_clock),
    .io_address(spriteMemories_30_io_address),
    .io_dataRead(spriteMemories_30_io_dataRead)
  );
  Memory_98 spriteMemories_31 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_31_clock),
    .io_address(spriteMemories_31_io_address),
    .io_dataRead(spriteMemories_31_io_dataRead)
  );
  Memory_99 spriteMemories_32 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_32_clock),
    .io_address(spriteMemories_32_io_address),
    .io_dataRead(spriteMemories_32_io_dataRead)
  );
  Memory_100 spriteMemories_33 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_33_clock),
    .io_address(spriteMemories_33_io_address),
    .io_dataRead(spriteMemories_33_io_dataRead)
  );
  Memory_101 spriteMemories_34 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_34_clock),
    .io_address(spriteMemories_34_io_address),
    .io_dataRead(spriteMemories_34_io_dataRead)
  );
  Memory_102 spriteMemories_35 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_35_clock),
    .io_address(spriteMemories_35_io_address),
    .io_dataRead(spriteMemories_35_io_dataRead)
  );
  Memory_103 spriteMemories_36 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_36_clock),
    .io_address(spriteMemories_36_io_address),
    .io_dataRead(spriteMemories_36_io_dataRead)
  );
  Memory_104 spriteMemories_37 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_37_clock),
    .io_address(spriteMemories_37_io_address),
    .io_dataRead(spriteMemories_37_io_dataRead)
  );
  Memory_105 spriteMemories_38 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_38_clock),
    .io_address(spriteMemories_38_io_address),
    .io_dataRead(spriteMemories_38_io_dataRead)
  );
  Memory_106 spriteMemories_39 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_39_clock),
    .io_address(spriteMemories_39_io_address),
    .io_dataRead(spriteMemories_39_io_dataRead)
  );
  Memory_107 spriteMemories_40 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_40_clock),
    .io_address(spriteMemories_40_io_address),
    .io_dataRead(spriteMemories_40_io_dataRead)
  );
  Memory_108 spriteMemories_41 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_41_clock),
    .io_address(spriteMemories_41_io_address),
    .io_dataRead(spriteMemories_41_io_dataRead)
  );
  Memory_109 spriteMemories_42 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_42_clock),
    .io_address(spriteMemories_42_io_address),
    .io_dataRead(spriteMemories_42_io_dataRead)
  );
  Memory_110 spriteMemories_43 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_43_clock),
    .io_address(spriteMemories_43_io_address),
    .io_dataRead(spriteMemories_43_io_dataRead)
  );
  Memory_111 spriteMemories_44 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_44_clock),
    .io_address(spriteMemories_44_io_address),
    .io_dataRead(spriteMemories_44_io_dataRead)
  );
  Memory_112 spriteMemories_45 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_45_clock),
    .io_address(spriteMemories_45_io_address),
    .io_dataRead(spriteMemories_45_io_dataRead)
  );
  Memory_113 spriteMemories_46 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_46_clock),
    .io_address(spriteMemories_46_io_address),
    .io_dataRead(spriteMemories_46_io_dataRead)
  );
  Memory_114 spriteMemories_47 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_47_clock),
    .io_address(spriteMemories_47_io_address),
    .io_dataRead(spriteMemories_47_io_dataRead)
  );
  Memory_115 spriteMemories_48 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_48_clock),
    .io_address(spriteMemories_48_io_address),
    .io_dataRead(spriteMemories_48_io_dataRead)
  );
  Memory_116 spriteMemories_49 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_49_clock),
    .io_address(spriteMemories_49_io_address),
    .io_dataRead(spriteMemories_49_io_dataRead)
  );
  Memory_117 spriteMemories_50 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_50_clock),
    .io_address(spriteMemories_50_io_address),
    .io_dataRead(spriteMemories_50_io_dataRead)
  );
  Memory_118 spriteMemories_51 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_51_clock),
    .io_address(spriteMemories_51_io_address),
    .io_dataRead(spriteMemories_51_io_dataRead)
  );
  Memory_119 spriteMemories_52 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_52_clock),
    .io_address(spriteMemories_52_io_address),
    .io_dataRead(spriteMemories_52_io_dataRead)
  );
  Memory_120 spriteMemories_53 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_53_clock),
    .io_address(spriteMemories_53_io_address),
    .io_dataRead(spriteMemories_53_io_dataRead)
  );
  Memory_121 spriteMemories_54 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_54_clock),
    .io_address(spriteMemories_54_io_address),
    .io_dataRead(spriteMemories_54_io_dataRead)
  );
  Memory_122 spriteMemories_55 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_55_clock),
    .io_address(spriteMemories_55_io_address),
    .io_dataRead(spriteMemories_55_io_dataRead)
  );
  Memory_123 spriteMemories_56 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_56_clock),
    .io_address(spriteMemories_56_io_address),
    .io_dataRead(spriteMemories_56_io_dataRead)
  );
  Memory_124 spriteMemories_57 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_57_clock),
    .io_address(spriteMemories_57_io_address),
    .io_dataRead(spriteMemories_57_io_dataRead)
  );
  Memory_125 spriteMemories_58 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_58_clock),
    .io_address(spriteMemories_58_io_address),
    .io_dataRead(spriteMemories_58_io_dataRead)
  );
  Memory_126 spriteMemories_59 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_59_clock),
    .io_address(spriteMemories_59_io_address),
    .io_dataRead(spriteMemories_59_io_dataRead)
  );
  Memory_127 spriteMemories_60 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_60_clock),
    .io_address(spriteMemories_60_io_address),
    .io_dataRead(spriteMemories_60_io_dataRead)
  );
  Memory_128 spriteMemories_61 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_61_clock),
    .io_address(spriteMemories_61_io_address),
    .io_dataRead(spriteMemories_61_io_dataRead)
  );
  Memory_129 spriteMemories_62 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_62_clock),
    .io_address(spriteMemories_62_io_address),
    .io_dataRead(spriteMemories_62_io_dataRead)
  );
  Memory_130 spriteMemories_63 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_63_clock),
    .io_address(spriteMemories_63_io_address),
    .io_dataRead(spriteMemories_63_io_dataRead)
  );
  MultiHotPriortyReductionTree multiHotPriortyReductionTree ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
    .io_dataInput_0(multiHotPriortyReductionTree_io_dataInput_0),
    .io_dataInput_1(multiHotPriortyReductionTree_io_dataInput_1),
    .io_dataInput_2(multiHotPriortyReductionTree_io_dataInput_2),
    .io_dataInput_3(multiHotPriortyReductionTree_io_dataInput_3),
    .io_dataInput_4(multiHotPriortyReductionTree_io_dataInput_4),
    .io_dataInput_5(multiHotPriortyReductionTree_io_dataInput_5),
    .io_dataInput_6(multiHotPriortyReductionTree_io_dataInput_6),
    .io_dataInput_7(multiHotPriortyReductionTree_io_dataInput_7),
    .io_dataInput_8(multiHotPriortyReductionTree_io_dataInput_8),
    .io_dataInput_9(multiHotPriortyReductionTree_io_dataInput_9),
    .io_dataInput_10(multiHotPriortyReductionTree_io_dataInput_10),
    .io_dataInput_11(multiHotPriortyReductionTree_io_dataInput_11),
    .io_dataInput_12(multiHotPriortyReductionTree_io_dataInput_12),
    .io_dataInput_13(multiHotPriortyReductionTree_io_dataInput_13),
    .io_dataInput_14(multiHotPriortyReductionTree_io_dataInput_14),
    .io_dataInput_15(multiHotPriortyReductionTree_io_dataInput_15),
    .io_dataInput_16(multiHotPriortyReductionTree_io_dataInput_16),
    .io_dataInput_17(multiHotPriortyReductionTree_io_dataInput_17),
    .io_dataInput_18(multiHotPriortyReductionTree_io_dataInput_18),
    .io_dataInput_19(multiHotPriortyReductionTree_io_dataInput_19),
    .io_dataInput_20(multiHotPriortyReductionTree_io_dataInput_20),
    .io_dataInput_21(multiHotPriortyReductionTree_io_dataInput_21),
    .io_dataInput_22(multiHotPriortyReductionTree_io_dataInput_22),
    .io_dataInput_23(multiHotPriortyReductionTree_io_dataInput_23),
    .io_dataInput_24(multiHotPriortyReductionTree_io_dataInput_24),
    .io_dataInput_25(multiHotPriortyReductionTree_io_dataInput_25),
    .io_dataInput_26(multiHotPriortyReductionTree_io_dataInput_26),
    .io_dataInput_27(multiHotPriortyReductionTree_io_dataInput_27),
    .io_dataInput_28(multiHotPriortyReductionTree_io_dataInput_28),
    .io_dataInput_29(multiHotPriortyReductionTree_io_dataInput_29),
    .io_dataInput_30(multiHotPriortyReductionTree_io_dataInput_30),
    .io_dataInput_31(multiHotPriortyReductionTree_io_dataInput_31),
    .io_dataInput_32(multiHotPriortyReductionTree_io_dataInput_32),
    .io_dataInput_33(multiHotPriortyReductionTree_io_dataInput_33),
    .io_dataInput_34(multiHotPriortyReductionTree_io_dataInput_34),
    .io_dataInput_35(multiHotPriortyReductionTree_io_dataInput_35),
    .io_dataInput_36(multiHotPriortyReductionTree_io_dataInput_36),
    .io_dataInput_37(multiHotPriortyReductionTree_io_dataInput_37),
    .io_dataInput_38(multiHotPriortyReductionTree_io_dataInput_38),
    .io_dataInput_39(multiHotPriortyReductionTree_io_dataInput_39),
    .io_dataInput_40(multiHotPriortyReductionTree_io_dataInput_40),
    .io_dataInput_41(multiHotPriortyReductionTree_io_dataInput_41),
    .io_dataInput_42(multiHotPriortyReductionTree_io_dataInput_42),
    .io_dataInput_43(multiHotPriortyReductionTree_io_dataInput_43),
    .io_dataInput_44(multiHotPriortyReductionTree_io_dataInput_44),
    .io_dataInput_45(multiHotPriortyReductionTree_io_dataInput_45),
    .io_dataInput_46(multiHotPriortyReductionTree_io_dataInput_46),
    .io_dataInput_47(multiHotPriortyReductionTree_io_dataInput_47),
    .io_dataInput_48(multiHotPriortyReductionTree_io_dataInput_48),
    .io_dataInput_49(multiHotPriortyReductionTree_io_dataInput_49),
    .io_dataInput_50(multiHotPriortyReductionTree_io_dataInput_50),
    .io_dataInput_51(multiHotPriortyReductionTree_io_dataInput_51),
    .io_dataInput_52(multiHotPriortyReductionTree_io_dataInput_52),
    .io_dataInput_53(multiHotPriortyReductionTree_io_dataInput_53),
    .io_dataInput_54(multiHotPriortyReductionTree_io_dataInput_54),
    .io_dataInput_55(multiHotPriortyReductionTree_io_dataInput_55),
    .io_dataInput_56(multiHotPriortyReductionTree_io_dataInput_56),
    .io_dataInput_57(multiHotPriortyReductionTree_io_dataInput_57),
    .io_dataInput_58(multiHotPriortyReductionTree_io_dataInput_58),
    .io_dataInput_59(multiHotPriortyReductionTree_io_dataInput_59),
    .io_dataInput_60(multiHotPriortyReductionTree_io_dataInput_60),
    .io_dataInput_61(multiHotPriortyReductionTree_io_dataInput_61),
    .io_dataInput_62(multiHotPriortyReductionTree_io_dataInput_62),
    .io_dataInput_63(multiHotPriortyReductionTree_io_dataInput_63),
    .io_selectInput_0(multiHotPriortyReductionTree_io_selectInput_0),
    .io_selectInput_1(multiHotPriortyReductionTree_io_selectInput_1),
    .io_selectInput_2(multiHotPriortyReductionTree_io_selectInput_2),
    .io_selectInput_3(multiHotPriortyReductionTree_io_selectInput_3),
    .io_selectInput_4(multiHotPriortyReductionTree_io_selectInput_4),
    .io_selectInput_5(multiHotPriortyReductionTree_io_selectInput_5),
    .io_selectInput_6(multiHotPriortyReductionTree_io_selectInput_6),
    .io_selectInput_7(multiHotPriortyReductionTree_io_selectInput_7),
    .io_selectInput_8(multiHotPriortyReductionTree_io_selectInput_8),
    .io_selectInput_9(multiHotPriortyReductionTree_io_selectInput_9),
    .io_selectInput_10(multiHotPriortyReductionTree_io_selectInput_10),
    .io_selectInput_11(multiHotPriortyReductionTree_io_selectInput_11),
    .io_selectInput_12(multiHotPriortyReductionTree_io_selectInput_12),
    .io_selectInput_13(multiHotPriortyReductionTree_io_selectInput_13),
    .io_selectInput_14(multiHotPriortyReductionTree_io_selectInput_14),
    .io_selectInput_15(multiHotPriortyReductionTree_io_selectInput_15),
    .io_selectInput_16(multiHotPriortyReductionTree_io_selectInput_16),
    .io_selectInput_17(multiHotPriortyReductionTree_io_selectInput_17),
    .io_selectInput_18(multiHotPriortyReductionTree_io_selectInput_18),
    .io_selectInput_19(multiHotPriortyReductionTree_io_selectInput_19),
    .io_selectInput_20(multiHotPriortyReductionTree_io_selectInput_20),
    .io_selectInput_21(multiHotPriortyReductionTree_io_selectInput_21),
    .io_selectInput_22(multiHotPriortyReductionTree_io_selectInput_22),
    .io_selectInput_23(multiHotPriortyReductionTree_io_selectInput_23),
    .io_selectInput_24(multiHotPriortyReductionTree_io_selectInput_24),
    .io_selectInput_25(multiHotPriortyReductionTree_io_selectInput_25),
    .io_selectInput_26(multiHotPriortyReductionTree_io_selectInput_26),
    .io_selectInput_27(multiHotPriortyReductionTree_io_selectInput_27),
    .io_selectInput_28(multiHotPriortyReductionTree_io_selectInput_28),
    .io_selectInput_29(multiHotPriortyReductionTree_io_selectInput_29),
    .io_selectInput_30(multiHotPriortyReductionTree_io_selectInput_30),
    .io_selectInput_31(multiHotPriortyReductionTree_io_selectInput_31),
    .io_selectInput_32(multiHotPriortyReductionTree_io_selectInput_32),
    .io_selectInput_33(multiHotPriortyReductionTree_io_selectInput_33),
    .io_selectInput_34(multiHotPriortyReductionTree_io_selectInput_34),
    .io_selectInput_35(multiHotPriortyReductionTree_io_selectInput_35),
    .io_selectInput_36(multiHotPriortyReductionTree_io_selectInput_36),
    .io_selectInput_37(multiHotPriortyReductionTree_io_selectInput_37),
    .io_selectInput_38(multiHotPriortyReductionTree_io_selectInput_38),
    .io_selectInput_39(multiHotPriortyReductionTree_io_selectInput_39),
    .io_selectInput_40(multiHotPriortyReductionTree_io_selectInput_40),
    .io_selectInput_41(multiHotPriortyReductionTree_io_selectInput_41),
    .io_selectInput_42(multiHotPriortyReductionTree_io_selectInput_42),
    .io_selectInput_43(multiHotPriortyReductionTree_io_selectInput_43),
    .io_selectInput_44(multiHotPriortyReductionTree_io_selectInput_44),
    .io_selectInput_45(multiHotPriortyReductionTree_io_selectInput_45),
    .io_selectInput_46(multiHotPriortyReductionTree_io_selectInput_46),
    .io_selectInput_47(multiHotPriortyReductionTree_io_selectInput_47),
    .io_selectInput_48(multiHotPriortyReductionTree_io_selectInput_48),
    .io_selectInput_49(multiHotPriortyReductionTree_io_selectInput_49),
    .io_selectInput_50(multiHotPriortyReductionTree_io_selectInput_50),
    .io_selectInput_51(multiHotPriortyReductionTree_io_selectInput_51),
    .io_selectInput_52(multiHotPriortyReductionTree_io_selectInput_52),
    .io_selectInput_53(multiHotPriortyReductionTree_io_selectInput_53),
    .io_selectInput_54(multiHotPriortyReductionTree_io_selectInput_54),
    .io_selectInput_55(multiHotPriortyReductionTree_io_selectInput_55),
    .io_selectInput_56(multiHotPriortyReductionTree_io_selectInput_56),
    .io_selectInput_57(multiHotPriortyReductionTree_io_selectInput_57),
    .io_selectInput_58(multiHotPriortyReductionTree_io_selectInput_58),
    .io_selectInput_59(multiHotPriortyReductionTree_io_selectInput_59),
    .io_selectInput_60(multiHotPriortyReductionTree_io_selectInput_60),
    .io_selectInput_61(multiHotPriortyReductionTree_io_selectInput_61),
    .io_selectInput_62(multiHotPriortyReductionTree_io_selectInput_62),
    .io_selectInput_63(multiHotPriortyReductionTree_io_selectInput_63),
    .io_dataOutput(multiHotPriortyReductionTree_io_dataOutput),
    .io_selectOutput(multiHotPriortyReductionTree_io_selectOutput)
  );
  assign io_newFrame = run & _GEN_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13 71:15]
  assign io_missingFrameError = missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 131:24]
  assign io_viewBoxOutOfRangeError = viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 133:29]
  assign io_vgaRed = io_vgaRed_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 349:13]
  assign io_vgaBlue = io_vgaBlue_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 351:14]
  assign io_vgaGreen = io_vgaGreen_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 350:15]
  assign io_Hsync = io_Hsync_pipeReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 94:12]
  assign io_Vsync = io_Vsync_pipeReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 95:12]
  assign backTileMemories_0_clock = clock;
  assign backTileMemories_0_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_1_clock = clock;
  assign backTileMemories_1_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_2_clock = clock;
  assign backTileMemories_2_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_3_clock = clock;
  assign backTileMemories_3_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_4_clock = clock;
  assign backTileMemories_4_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_5_clock = clock;
  assign backTileMemories_5_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_6_clock = clock;
  assign backTileMemories_6_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_7_clock = clock;
  assign backTileMemories_7_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_8_clock = clock;
  assign backTileMemories_8_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_9_clock = clock;
  assign backTileMemories_9_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_10_clock = clock;
  assign backTileMemories_10_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_11_clock = clock;
  assign backTileMemories_11_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_12_clock = clock;
  assign backTileMemories_12_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_13_clock = clock;
  assign backTileMemories_13_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_14_clock = clock;
  assign backTileMemories_14_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_15_clock = clock;
  assign backTileMemories_15_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_16_clock = clock;
  assign backTileMemories_16_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_17_clock = clock;
  assign backTileMemories_17_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_18_clock = clock;
  assign backTileMemories_18_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_19_clock = clock;
  assign backTileMemories_19_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_20_clock = clock;
  assign backTileMemories_20_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_21_clock = clock;
  assign backTileMemories_21_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_22_clock = clock;
  assign backTileMemories_22_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_23_clock = clock;
  assign backTileMemories_23_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_24_clock = clock;
  assign backTileMemories_24_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_25_clock = clock;
  assign backTileMemories_25_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_26_clock = clock;
  assign backTileMemories_26_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_27_clock = clock;
  assign backTileMemories_27_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_28_clock = clock;
  assign backTileMemories_28_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_29_clock = clock;
  assign backTileMemories_29_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_30_clock = clock;
  assign backTileMemories_30_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_31_clock = clock;
  assign backTileMemories_31_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_32_clock = clock;
  assign backTileMemories_32_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_33_clock = clock;
  assign backTileMemories_33_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_34_clock = clock;
  assign backTileMemories_34_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_35_clock = clock;
  assign backTileMemories_35_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_36_clock = clock;
  assign backTileMemories_36_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_37_clock = clock;
  assign backTileMemories_37_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_38_clock = clock;
  assign backTileMemories_38_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_39_clock = clock;
  assign backTileMemories_39_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_40_clock = clock;
  assign backTileMemories_40_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_41_clock = clock;
  assign backTileMemories_41_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_42_clock = clock;
  assign backTileMemories_42_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_43_clock = clock;
  assign backTileMemories_43_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_44_clock = clock;
  assign backTileMemories_44_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_45_clock = clock;
  assign backTileMemories_45_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_46_clock = clock;
  assign backTileMemories_46_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_47_clock = clock;
  assign backTileMemories_47_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_48_clock = clock;
  assign backTileMemories_48_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_49_clock = clock;
  assign backTileMemories_49_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_50_clock = clock;
  assign backTileMemories_50_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_51_clock = clock;
  assign backTileMemories_51_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_52_clock = clock;
  assign backTileMemories_52_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_53_clock = clock;
  assign backTileMemories_53_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_54_clock = clock;
  assign backTileMemories_54_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_55_clock = clock;
  assign backTileMemories_55_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_56_clock = clock;
  assign backTileMemories_56_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_57_clock = clock;
  assign backTileMemories_57_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_58_clock = clock;
  assign backTileMemories_58_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_59_clock = clock;
  assign backTileMemories_59_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_60_clock = clock;
  assign backTileMemories_60_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_61_clock = clock;
  assign backTileMemories_61_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_62_clock = clock;
  assign backTileMemories_62_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_63_clock = clock;
  assign backTileMemories_63_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backBufferMemory_clock = clock;
  assign backBufferMemory_io_address = _backBufferMemory_io_address_T_5[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:31]
  assign backBufferMemory_io_writeEnable = copyEnabledReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 228:35]
  assign backBufferMemory_io_dataWrite = backBufferShadowMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 229:33]
  assign backBufferShadowMemory_clock = clock;
  assign backBufferShadowMemory_io_address = restoreEnabled ? backBufferShadowMemory_io_address_REG :
    _backBufferShadowMemory_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:43]
  assign backBufferShadowMemory_io_writeEnable = restoreEnabled & backBufferShadowMemory_io_writeEnable_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:47]
  assign backBufferShadowMemory_io_dataWrite = restoreEnabled ? backBufferRestoreMemory_io_dataRead : 6'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 224:45]
  assign backBufferRestoreMemory_clock = clock;
  assign backBufferRestoreMemory_io_address = backMemoryRestoreCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 216:65]
  assign spriteMemories_0_clock = clock;
  assign spriteMemories_0_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_1_clock = clock;
  assign spriteMemories_1_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_2_clock = clock;
  assign spriteMemories_2_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_3_clock = clock;
  assign spriteMemories_3_io_address = _spriteMemories_3_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_4_clock = clock;
  assign spriteMemories_4_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_5_clock = clock;
  assign spriteMemories_5_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_6_clock = clock;
  assign spriteMemories_6_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_7_clock = clock;
  assign spriteMemories_7_io_address = _spriteMemories_7_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_8_clock = clock;
  assign spriteMemories_8_io_address = _spriteMemories_8_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_9_clock = clock;
  assign spriteMemories_9_io_address = _spriteMemories_9_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_10_clock = clock;
  assign spriteMemories_10_io_address = _spriteMemories_10_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_11_clock = clock;
  assign spriteMemories_11_io_address = _spriteMemories_11_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_12_clock = clock;
  assign spriteMemories_12_io_address = _spriteMemories_12_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_13_clock = clock;
  assign spriteMemories_13_io_address = _spriteMemories_13_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_14_clock = clock;
  assign spriteMemories_14_io_address = _spriteMemories_14_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_15_clock = clock;
  assign spriteMemories_15_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_16_clock = clock;
  assign spriteMemories_16_io_address = _spriteMemories_16_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_17_clock = clock;
  assign spriteMemories_17_io_address = _spriteMemories_17_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_18_clock = clock;
  assign spriteMemories_18_io_address = _spriteMemories_18_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_19_clock = clock;
  assign spriteMemories_19_io_address = _spriteMemories_19_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_20_clock = clock;
  assign spriteMemories_20_io_address = _spriteMemories_20_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_21_clock = clock;
  assign spriteMemories_21_io_address = _spriteMemories_21_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_22_clock = clock;
  assign spriteMemories_22_io_address = _spriteMemories_22_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_23_clock = clock;
  assign spriteMemories_23_io_address = _spriteMemories_23_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_24_clock = clock;
  assign spriteMemories_24_io_address = _spriteMemories_24_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_25_clock = clock;
  assign spriteMemories_25_io_address = _spriteMemories_25_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_26_clock = clock;
  assign spriteMemories_26_io_address = _spriteMemories_26_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_27_clock = clock;
  assign spriteMemories_27_io_address = _spriteMemories_27_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_28_clock = clock;
  assign spriteMemories_28_io_address = _spriteMemories_28_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_29_clock = clock;
  assign spriteMemories_29_io_address = _spriteMemories_29_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_30_clock = clock;
  assign spriteMemories_30_io_address = _spriteMemories_30_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_31_clock = clock;
  assign spriteMemories_31_io_address = _spriteMemories_31_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_32_clock = clock;
  assign spriteMemories_32_io_address = _spriteMemories_32_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_33_clock = clock;
  assign spriteMemories_33_io_address = _spriteMemories_33_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_34_clock = clock;
  assign spriteMemories_34_io_address = _spriteMemories_34_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_35_clock = clock;
  assign spriteMemories_35_io_address = _spriteMemories_35_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_36_clock = clock;
  assign spriteMemories_36_io_address = _spriteMemories_36_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_37_clock = clock;
  assign spriteMemories_37_io_address = _spriteMemories_37_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_38_clock = clock;
  assign spriteMemories_38_io_address = _spriteMemories_38_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_39_clock = clock;
  assign spriteMemories_39_io_address = _spriteMemories_39_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_40_clock = clock;
  assign spriteMemories_40_io_address = _spriteMemories_40_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_41_clock = clock;
  assign spriteMemories_41_io_address = _spriteMemories_41_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_42_clock = clock;
  assign spriteMemories_42_io_address = _spriteMemories_42_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_43_clock = clock;
  assign spriteMemories_43_io_address = _spriteMemories_43_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_44_clock = clock;
  assign spriteMemories_44_io_address = _spriteMemories_44_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_45_clock = clock;
  assign spriteMemories_45_io_address = _spriteMemories_45_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_46_clock = clock;
  assign spriteMemories_46_io_address = _spriteMemories_46_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_47_clock = clock;
  assign spriteMemories_47_io_address = _spriteMemories_47_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_48_clock = clock;
  assign spriteMemories_48_io_address = _spriteMemories_48_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_49_clock = clock;
  assign spriteMemories_49_io_address = _spriteMemories_49_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_50_clock = clock;
  assign spriteMemories_50_io_address = _spriteMemories_50_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_51_clock = clock;
  assign spriteMemories_51_io_address = _spriteMemories_51_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_52_clock = clock;
  assign spriteMemories_52_io_address = _spriteMemories_52_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_53_clock = clock;
  assign spriteMemories_53_io_address = _spriteMemories_53_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_54_clock = clock;
  assign spriteMemories_54_io_address = _spriteMemories_54_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_55_clock = clock;
  assign spriteMemories_55_io_address = _spriteMemories_55_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_56_clock = clock;
  assign spriteMemories_56_io_address = _spriteMemories_56_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_57_clock = clock;
  assign spriteMemories_57_io_address = _spriteMemories_57_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_58_clock = clock;
  assign spriteMemories_58_io_address = _spriteMemories_58_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_59_clock = clock;
  assign spriteMemories_59_io_address = _spriteMemories_59_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_60_clock = clock;
  assign spriteMemories_60_io_address = _spriteMemories_60_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_61_clock = clock;
  assign spriteMemories_61_io_address = _spriteMemories_61_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_62_clock = clock;
  assign spriteMemories_62_io_address = _spriteMemories_62_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_63_clock = clock;
  assign spriteMemories_63_io_address = _spriteMemories_63_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign multiHotPriortyReductionTree_io_dataInput_0 = multiHotPriortyReductionTree_io_dataInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_1 = multiHotPriortyReductionTree_io_dataInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_2 = multiHotPriortyReductionTree_io_dataInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_3 = multiHotPriortyReductionTree_io_dataInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_4 = multiHotPriortyReductionTree_io_dataInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_5 = multiHotPriortyReductionTree_io_dataInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_6 = multiHotPriortyReductionTree_io_dataInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_7 = multiHotPriortyReductionTree_io_dataInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_8 = multiHotPriortyReductionTree_io_dataInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_9 = multiHotPriortyReductionTree_io_dataInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_10 = multiHotPriortyReductionTree_io_dataInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_11 = multiHotPriortyReductionTree_io_dataInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_12 = multiHotPriortyReductionTree_io_dataInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_13 = multiHotPriortyReductionTree_io_dataInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_14 = multiHotPriortyReductionTree_io_dataInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_15 = multiHotPriortyReductionTree_io_dataInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_16 = multiHotPriortyReductionTree_io_dataInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_17 = multiHotPriortyReductionTree_io_dataInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_18 = multiHotPriortyReductionTree_io_dataInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_19 = multiHotPriortyReductionTree_io_dataInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_20 = multiHotPriortyReductionTree_io_dataInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_21 = multiHotPriortyReductionTree_io_dataInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_22 = multiHotPriortyReductionTree_io_dataInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_23 = multiHotPriortyReductionTree_io_dataInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_24 = multiHotPriortyReductionTree_io_dataInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_25 = multiHotPriortyReductionTree_io_dataInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_26 = multiHotPriortyReductionTree_io_dataInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_27 = multiHotPriortyReductionTree_io_dataInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_28 = multiHotPriortyReductionTree_io_dataInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_29 = multiHotPriortyReductionTree_io_dataInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_30 = multiHotPriortyReductionTree_io_dataInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_31 = multiHotPriortyReductionTree_io_dataInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_32 = multiHotPriortyReductionTree_io_dataInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_33 = multiHotPriortyReductionTree_io_dataInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_34 = multiHotPriortyReductionTree_io_dataInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_35 = multiHotPriortyReductionTree_io_dataInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_36 = multiHotPriortyReductionTree_io_dataInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_37 = multiHotPriortyReductionTree_io_dataInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_38 = multiHotPriortyReductionTree_io_dataInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_39 = multiHotPriortyReductionTree_io_dataInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_40 = multiHotPriortyReductionTree_io_dataInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_41 = multiHotPriortyReductionTree_io_dataInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_42 = multiHotPriortyReductionTree_io_dataInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_43 = multiHotPriortyReductionTree_io_dataInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_44 = multiHotPriortyReductionTree_io_dataInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_45 = multiHotPriortyReductionTree_io_dataInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_46 = multiHotPriortyReductionTree_io_dataInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_47 = multiHotPriortyReductionTree_io_dataInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_48 = multiHotPriortyReductionTree_io_dataInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_49 = multiHotPriortyReductionTree_io_dataInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_50 = multiHotPriortyReductionTree_io_dataInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_51 = multiHotPriortyReductionTree_io_dataInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_52 = multiHotPriortyReductionTree_io_dataInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_53 = multiHotPriortyReductionTree_io_dataInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_54 = multiHotPriortyReductionTree_io_dataInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_55 = multiHotPriortyReductionTree_io_dataInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_56 = multiHotPriortyReductionTree_io_dataInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_57 = multiHotPriortyReductionTree_io_dataInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_58 = multiHotPriortyReductionTree_io_dataInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_59 = multiHotPriortyReductionTree_io_dataInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_60 = multiHotPriortyReductionTree_io_dataInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_61 = multiHotPriortyReductionTree_io_dataInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_62 = multiHotPriortyReductionTree_io_dataInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_63 = multiHotPriortyReductionTree_io_dataInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_selectInput_0 = multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_1 = multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_2 = multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_3 = multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_4 = multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_5 = multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_6 = multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_7 = multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_8 = multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_9 = multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_10 = multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_11 = multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_12 = multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_13 = multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_14 = multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_15 = multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_16 = multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_17 = multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_18 = multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_19 = multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_20 = multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_21 = multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_22 = multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_23 = multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_24 = multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_25 = multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_26 = multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_27 = multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_28 = multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_29 = multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_30 = multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_31 = multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_32 = multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_32_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_33 = multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_33_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_34 = multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_34_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_35 = multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_35_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_36 = multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_36_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_37 = multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_37_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_38 = multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_38_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_39 = multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_39_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_40 = multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_40_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_41 = multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_41_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_42 = multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_42_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_43 = multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_43_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_44 = multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_44_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_45 = multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_45_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_46 = multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_46_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_47 = multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_47_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_48 = multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_48_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_49 = multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_49_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_50 = multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_50_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_51 = multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_51_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_52 = multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_52_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_53 = multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_53_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_54 = multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_54_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_55 = multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_55_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_56 = multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_56_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_57 = multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_57_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_58 = multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_58_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_59 = multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_59_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_60 = multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_60_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_61 = multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_61_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_62 = multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_62_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_63 = multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_63_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
      ScaleCounterReg <= 2'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        ScaleCounterReg <= 2'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 75:23]
      end else begin
        ScaleCounterReg <= _ScaleCounterReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 88:23]
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
      CounterXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        if (CounterXReg == 10'h31f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129]
          CounterXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 77:21]
        end else begin
          CounterXReg <= _CounterXReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 85:21]
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
      CounterYReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        if (CounterXReg == 10'h31f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129]
          CounterYReg <= _GEN_0;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
      backMemoryRestoreCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
    end else if (restoreEnabled) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:70]
      backMemoryRestoreCounter <= _backMemoryRestoreCounter_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 206:30]
    end
    io_Hsync_pipeReg_0 <= io_Hsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_1 <= io_Hsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_2 <= io_Hsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_3 <= ~Hsync; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 94:27]
    io_Vsync_pipeReg_0 <= io_Vsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_1 <= io_Vsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_2 <= io_Vsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_3 <= ~Vsync; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 95:27]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
      frameClockCount <= 21'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
    end else if (frameClockCount == 21'h19a27f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 105:25]
      frameClockCount <= 21'h0;
    end else begin
      frameClockCount <= _frameClockCount_T_2;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_3 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_3 <= io_spriteXPosition_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_7 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_7 <= io_spriteXPosition_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_8 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_8 <= io_spriteXPosition_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_9 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_9 <= io_spriteXPosition_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_10 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_10 <= io_spriteXPosition_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_11 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_11 <= io_spriteXPosition_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_12 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_12 <= io_spriteXPosition_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_13 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_13 <= io_spriteXPosition_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_14 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_14 <= io_spriteXPosition_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_16 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_16 <= io_spriteXPosition_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_17 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_17 <= io_spriteXPosition_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_18 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_18 <= io_spriteXPosition_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_19 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_19 <= io_spriteXPosition_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_20 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_20 <= io_spriteXPosition_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_21 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_21 <= io_spriteXPosition_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_22 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_22 <= io_spriteXPosition_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_23 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_23 <= io_spriteXPosition_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_24 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_24 <= io_spriteXPosition_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_25 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_25 <= io_spriteXPosition_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_26 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_26 <= io_spriteXPosition_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_27 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_27 <= io_spriteXPosition_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_28 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_28 <= io_spriteXPosition_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_29 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_29 <= io_spriteXPosition_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_30 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_30 <= io_spriteXPosition_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_31 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_31 <= io_spriteXPosition_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_32 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_32 <= io_spriteXPosition_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_33 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_33 <= io_spriteXPosition_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_34 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_34 <= io_spriteXPosition_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_35 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_35 <= io_spriteXPosition_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_36 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_36 <= io_spriteXPosition_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_37 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_37 <= io_spriteXPosition_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_38 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_38 <= io_spriteXPosition_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_39 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_39 <= io_spriteXPosition_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_40 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_40 <= io_spriteXPosition_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_41 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_41 <= io_spriteXPosition_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_42 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_42 <= io_spriteXPosition_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_43 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_43 <= io_spriteXPosition_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_44 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_44 <= io_spriteXPosition_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_45 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_45 <= io_spriteXPosition_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_46 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_46 <= io_spriteXPosition_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_47 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_47 <= io_spriteXPosition_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_48 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_48 <= io_spriteXPosition_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_49 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_49 <= io_spriteXPosition_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_50 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_50 <= io_spriteXPosition_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_51 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_51 <= io_spriteXPosition_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_52 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_52 <= io_spriteXPosition_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_53 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_53 <= io_spriteXPosition_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_54 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_54 <= io_spriteXPosition_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_55 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_55 <= io_spriteXPosition_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_56 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_56 <= io_spriteXPosition_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_57 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_57 <= io_spriteXPosition_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_58 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_58 <= io_spriteXPosition_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_59 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_59 <= io_spriteXPosition_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_60 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_60 <= io_spriteXPosition_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_61 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_61 <= io_spriteXPosition_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_62 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_62 <= io_spriteXPosition_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_63 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_63 <= io_spriteXPosition_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_3 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_3 <= io_spriteYPosition_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_7 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_7 <= io_spriteYPosition_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_8 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_8 <= io_spriteYPosition_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_9 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_9 <= io_spriteYPosition_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_10 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_10 <= io_spriteYPosition_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_11 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_11 <= io_spriteYPosition_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_12 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_12 <= io_spriteYPosition_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_13 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_13 <= io_spriteYPosition_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_14 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_14 <= io_spriteYPosition_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_16 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_16 <= io_spriteYPosition_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_17 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_17 <= io_spriteYPosition_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_18 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_18 <= io_spriteYPosition_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_19 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_19 <= io_spriteYPosition_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_20 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_20 <= io_spriteYPosition_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_21 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_21 <= io_spriteYPosition_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_22 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_22 <= io_spriteYPosition_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_23 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_23 <= io_spriteYPosition_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_24 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_24 <= io_spriteYPosition_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_25 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_25 <= io_spriteYPosition_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_26 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_26 <= io_spriteYPosition_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_27 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_27 <= io_spriteYPosition_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_28 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_28 <= io_spriteYPosition_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_29 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_29 <= io_spriteYPosition_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_30 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_30 <= io_spriteYPosition_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_31 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_31 <= io_spriteYPosition_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_32 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_32 <= io_spriteYPosition_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_33 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_33 <= io_spriteYPosition_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_34 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_34 <= io_spriteYPosition_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_35 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_35 <= io_spriteYPosition_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_36 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_36 <= io_spriteYPosition_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_37 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_37 <= io_spriteYPosition_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_38 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_38 <= io_spriteYPosition_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_39 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_39 <= io_spriteYPosition_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_40 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_40 <= io_spriteYPosition_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_41 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_41 <= io_spriteYPosition_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_42 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_42 <= io_spriteYPosition_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_43 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_43 <= io_spriteYPosition_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_44 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_44 <= io_spriteYPosition_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_45 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_45 <= io_spriteYPosition_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_46 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_46 <= io_spriteYPosition_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_47 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_47 <= io_spriteYPosition_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_48 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_48 <= io_spriteYPosition_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_49 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_49 <= io_spriteYPosition_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_50 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_50 <= io_spriteYPosition_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_51 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_51 <= io_spriteYPosition_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_52 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_52 <= io_spriteYPosition_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_53 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_53 <= io_spriteYPosition_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_54 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_54 <= io_spriteYPosition_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_55 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_55 <= io_spriteYPosition_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_56 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_56 <= io_spriteYPosition_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_57 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_57 <= io_spriteYPosition_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_58 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_58 <= io_spriteYPosition_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_59 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_59 <= io_spriteYPosition_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_60 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_60 <= io_spriteYPosition_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_61 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_61 <= io_spriteYPosition_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_62 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_62 <= io_spriteYPosition_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_63 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_63 <= io_spriteYPosition_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    spriteVisibleReg_0 <= reset | _GEN_141; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_1 <= reset | _GEN_142; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_2 <= reset | _GEN_143; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_3 <= reset | _GEN_144; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_4 <= reset | _GEN_145; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_5 <= reset | _GEN_146; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_6 <= reset | _GEN_147; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_7 <= reset | _GEN_148; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_8 <= reset | _GEN_149; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_9 <= reset | _GEN_150; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_10 <= reset | _GEN_151; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_11 <= reset | _GEN_152; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_12 <= reset | _GEN_153; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_13 <= reset | _GEN_154; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_14 <= reset | _GEN_155; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_15 <= reset | _GEN_156; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_16 <= reset | _GEN_157; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_17 <= reset | _GEN_158; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_18 <= reset | _GEN_159; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_19 <= reset | _GEN_160; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_20 <= reset | _GEN_161; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_21 <= reset | _GEN_162; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_22 <= reset | _GEN_163; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_23 <= reset | _GEN_164; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_24 <= reset | _GEN_165; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_25 <= reset | _GEN_166; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_26 <= reset | _GEN_167; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_27 <= reset | _GEN_168; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_28 <= reset | _GEN_169; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_29 <= reset | _GEN_170; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_30 <= reset | _GEN_171; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_31 <= reset | _GEN_172; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_32 <= reset | _GEN_173; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_33 <= reset | _GEN_174; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_34 <= reset | _GEN_175; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_35 <= reset | _GEN_176; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_36 <= reset | _GEN_177; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_37 <= reset | _GEN_178; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_38 <= reset | _GEN_179; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_39 <= reset | _GEN_180; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_40 <= reset | _GEN_181; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_41 <= reset | _GEN_182; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_42 <= reset | _GEN_183; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_43 <= reset | _GEN_184; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_44 <= reset | _GEN_185; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_45 <= reset | _GEN_186; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_46 <= reset | _GEN_187; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_47 <= reset | _GEN_188; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_48 <= reset | _GEN_189; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_49 <= reset | _GEN_190; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_50 <= reset | _GEN_191; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_51 <= reset | _GEN_192; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_52 <= reset | _GEN_193; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_53 <= reset | _GEN_194; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_54 <= reset | _GEN_195; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_55 <= reset | _GEN_196; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_56 <= reset | _GEN_197; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_57 <= reset | _GEN_198; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_58 <= reset | _GEN_199; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_59 <= reset | _GEN_200; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_60 <= reset | _GEN_201; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_61 <= reset | _GEN_202; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_62 <= reset | _GEN_203; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_63 <= reset | _GEN_204; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_16 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_16 <= io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_17 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_17 <= io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_18 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_18 <= io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_19 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_19 <= io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_20 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_20 <= io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_21 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_21 <= io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_22 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_22 <= io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_23 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_23 <= io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_24 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_24 <= io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_25 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_25 <= io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_26 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_26 <= io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_27 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_27 <= io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_28 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_28 <= io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_29 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_29 <= io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_30 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_30 <= io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_31 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_31 <= io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_32 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_32 <= io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_33 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_33 <= io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_34 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_34 <= io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_35 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_35 <= io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_36 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_36 <= io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_37 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_37 <= io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_38 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_38 <= io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_39 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_39 <= io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_40 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_40 <= io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_41 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_41 <= io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_42 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_42 <= io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_43 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_43 <= io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_44 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_44 <= io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_45 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_45 <= io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_58 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_58 <= io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_59 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_59 <= io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_60 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
      spriteScaleUpHorizontalReg_60 <= io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 119:45]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_16 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_16 <= io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_17 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_17 <= io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_18 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_18 <= io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_19 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_19 <= io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_20 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_20 <= io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_21 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_21 <= io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_22 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_22 <= io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_23 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_23 <= io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_24 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_24 <= io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_25 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_25 <= io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_26 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_26 <= io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_27 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_27 <= io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_28 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_28 <= io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_29 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_29 <= io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_30 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_30 <= io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_31 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_31 <= io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_32 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_32 <= io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_33 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_33 <= io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_34 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_34 <= io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_35 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_35 <= io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_36 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_36 <= io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_37 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_37 <= io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_38 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_38 <= io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_39 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_39 <= io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_40 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_40 <= io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_41 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_41 <= io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_42 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_42 <= io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_43 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_43 <= io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_44 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_44 <= io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_45 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_45 <= io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_58 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_58 <= io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_59 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_59 <= io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_60 <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
      spriteScaleUpVerticalReg_60 <= io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 121:43]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
      viewBoxXReg <= io_viewBoxX; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
      viewBoxYReg <= 9'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
      viewBoxYReg <= io_viewBoxY; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
      missingFrameErrorReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
    end else begin
      missingFrameErrorReg <= _GEN_594;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
      viewBoxOutOfRangeErrorReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
    end else begin
      viewBoxOutOfRangeErrorReg <= _GEN_591;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
      newFrameStikyReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
    end else if (REG) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:37]
      newFrameStikyReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 152:22]
    end else begin
      newFrameStikyReg <= _GEN_592;
    end
    REG <= io_frameUpdateDone; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:16]
    backTileMemoryDataRead_0_REG <= backTileMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_1_REG <= backTileMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_2_REG <= backTileMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_3_REG <= backTileMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_4_REG <= backTileMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_5_REG <= backTileMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_6_REG <= backTileMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_7_REG <= backTileMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_8_REG <= backTileMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_9_REG <= backTileMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_10_REG <= backTileMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_11_REG <= backTileMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_12_REG <= backTileMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_13_REG <= backTileMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_14_REG <= backTileMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_15_REG <= backTileMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_16_REG <= backTileMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_17_REG <= backTileMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_18_REG <= backTileMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_19_REG <= backTileMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_20_REG <= backTileMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_21_REG <= backTileMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_22_REG <= backTileMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_23_REG <= backTileMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_24_REG <= backTileMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_25_REG <= backTileMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_26_REG <= backTileMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_27_REG <= backTileMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_28_REG <= backTileMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_29_REG <= backTileMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_30_REG <= backTileMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_31_REG <= backTileMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_32_REG <= backTileMemories_32_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_33_REG <= backTileMemories_33_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_34_REG <= backTileMemories_34_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_35_REG <= backTileMemories_35_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_36_REG <= backTileMemories_36_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_37_REG <= backTileMemories_37_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_38_REG <= backTileMemories_38_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_39_REG <= backTileMemories_39_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_40_REG <= backTileMemories_40_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_41_REG <= backTileMemories_41_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_42_REG <= backTileMemories_42_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_43_REG <= backTileMemories_43_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_44_REG <= backTileMemories_44_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_45_REG <= backTileMemories_45_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_46_REG <= backTileMemories_46_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_47_REG <= backTileMemories_47_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_48_REG <= backTileMemories_48_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_49_REG <= backTileMemories_49_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_50_REG <= backTileMemories_50_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_51_REG <= backTileMemories_51_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_52_REG <= backTileMemories_52_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_53_REG <= backTileMemories_53_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_54_REG <= backTileMemories_54_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_55_REG <= backTileMemories_55_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_56_REG <= backTileMemories_56_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_57_REG <= backTileMemories_57_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_58_REG <= backTileMemories_58_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_59_REG <= backTileMemories_59_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_60_REG <= backTileMemories_60_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_61_REG <= backTileMemories_61_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_62_REG <= backTileMemories_62_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_63_REG <= backTileMemories_63_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
      backMemoryCopyCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
    end else if (preDisplayArea) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23]
      if (backMemoryCopyCounter < 12'h800) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 187:66]
        backMemoryCopyCounter <= _backMemoryCopyCounter_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 188:29]
      end
    end else begin
      backMemoryCopyCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 197:27]
    end
    copyEnabledReg <= preDisplayArea & _T_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23 198:17]
    backBufferShadowMemory_io_address_REG <= backMemoryRestoreCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:92]
    backBufferShadowMemory_io_writeEnable_REG <= backMemoryRestoreCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:33]
    backBufferMemory_io_address_REG <= backMemoryCopyCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:83]
    fullBackgroundColor_REG <= backBufferMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:56]
    if (fullBackgroundColor[6]) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 244:25]
      pixelColorBack <= 6'h0;
    end else begin
      pixelColorBack <= fullBackgroundColor[5:0];
    end
    multiHotPriortyReductionTree_io_dataInput_0_REG <= spriteMemories_0_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1 <= spriteVisibleReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_0_REG <= spriteMemories_0_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_1_REG <= spriteMemories_1_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1 <= spriteVisibleReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_1_REG <= spriteMemories_1_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_2_REG <= spriteMemories_2_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1 <= spriteVisibleReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_2_REG <= spriteMemories_2_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_3_REG <= spriteMemories_3_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1 <= spriteVisibleReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1 <= inSpriteHorizontal_3 & inSpriteVertical_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_3_REG <= spriteMemories_3_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_4_REG <= spriteMemories_4_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1 <= spriteVisibleReg_4; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_4_REG <= spriteMemories_4_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_5_REG <= spriteMemories_5_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1 <= spriteVisibleReg_5; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_5_REG <= spriteMemories_5_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_6_REG <= spriteMemories_6_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1 <= spriteVisibleReg_6; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_6_REG <= spriteMemories_6_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_7_REG <= spriteMemories_7_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1 <= spriteVisibleReg_7; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1 <= inSpriteHorizontal_7 & inSpriteVertical_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_7_REG <= spriteMemories_7_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_8_REG <= spriteMemories_8_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1 <= spriteVisibleReg_8; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1 <= inSpriteHorizontal_8 & inSpriteVertical_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_8_REG <= spriteMemories_8_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_9_REG <= spriteMemories_9_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1 <= spriteVisibleReg_9; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1 <= inSpriteHorizontal_9 & inSpriteVertical_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_9_REG <= spriteMemories_9_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_10_REG <= spriteMemories_10_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1 <= spriteVisibleReg_10; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1 <= inSpriteHorizontal_10 & inSpriteVertical_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_10_REG <= spriteMemories_10_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_11_REG <= spriteMemories_11_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1 <= spriteVisibleReg_11; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1 <= inSpriteHorizontal_11 & inSpriteVertical_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_11_REG <= spriteMemories_11_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_12_REG <= spriteMemories_12_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1 <= spriteVisibleReg_12; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1 <= inSpriteHorizontal_12 & inSpriteVertical_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_12_REG <= spriteMemories_12_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_13_REG <= spriteMemories_13_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1 <= spriteVisibleReg_13; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1 <= inSpriteHorizontal_13 & inSpriteVertical_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_13_REG <= spriteMemories_13_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_14_REG <= spriteMemories_14_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1 <= spriteVisibleReg_14; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1 <= inSpriteHorizontal_14 & inSpriteVertical_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_14_REG <= spriteMemories_14_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_15_REG <= spriteMemories_15_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1 <= spriteVisibleReg_15; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_15_REG <= spriteMemories_15_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_16_REG <= spriteMemories_16_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1 <= spriteVisibleReg_16; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1 <= inSpriteHorizontal_16 & inSpriteVertical_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_16_REG <= spriteMemories_16_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_17_REG <= spriteMemories_17_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1 <= spriteVisibleReg_17; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1 <= inSpriteHorizontal_17 & inSpriteVertical_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_17_REG <= spriteMemories_17_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_18_REG <= spriteMemories_18_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1 <= spriteVisibleReg_18; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1 <= inSpriteHorizontal_18 & inSpriteVertical_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_18_REG <= spriteMemories_18_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_19_REG <= spriteMemories_19_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1 <= spriteVisibleReg_19; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1 <= inSpriteHorizontal_19 & inSpriteVertical_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_19_REG <= spriteMemories_19_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_20_REG <= spriteMemories_20_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1 <= spriteVisibleReg_20; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1 <= inSpriteHorizontal_20 & inSpriteVertical_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_20_REG <= spriteMemories_20_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_21_REG <= spriteMemories_21_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1 <= spriteVisibleReg_21; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1 <= inSpriteHorizontal_21 & inSpriteVertical_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_21_REG <= spriteMemories_21_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_22_REG <= spriteMemories_22_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1 <= spriteVisibleReg_22; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1 <= inSpriteHorizontal_22 & inSpriteVertical_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_22_REG <= spriteMemories_22_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_23_REG <= spriteMemories_23_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1 <= spriteVisibleReg_23; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1 <= inSpriteHorizontal_23 & inSpriteVertical_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_23_REG <= spriteMemories_23_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_24_REG <= spriteMemories_24_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1 <= spriteVisibleReg_24; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1 <= inSpriteHorizontal_24 & inSpriteVertical_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_24_REG <= spriteMemories_24_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_25_REG <= spriteMemories_25_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1 <= spriteVisibleReg_25; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1 <= inSpriteHorizontal_25 & inSpriteVertical_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_25_REG <= spriteMemories_25_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_26_REG <= spriteMemories_26_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1 <= spriteVisibleReg_26; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1 <= inSpriteHorizontal_26 & inSpriteVertical_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_26_REG <= spriteMemories_26_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_27_REG <= spriteMemories_27_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1 <= spriteVisibleReg_27; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1 <= inSpriteHorizontal_27 & inSpriteVertical_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_27_REG <= spriteMemories_27_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_28_REG <= spriteMemories_28_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1 <= spriteVisibleReg_28; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1 <= inSpriteHorizontal_28 & inSpriteVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_28_REG <= spriteMemories_28_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_29_REG <= spriteMemories_29_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1 <= spriteVisibleReg_29; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1 <= inSpriteHorizontal_29 & inSpriteVertical_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_29_REG <= spriteMemories_29_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_30_REG <= spriteMemories_30_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1 <= spriteVisibleReg_30; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1 <= inSpriteHorizontal_30 & inSpriteVertical_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_30_REG <= spriteMemories_30_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_31_REG <= spriteMemories_31_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1 <= spriteVisibleReg_31; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1 <= inSpriteHorizontal_31 & inSpriteVertical_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_31_REG <= spriteMemories_31_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_32_REG <= spriteMemories_32_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1 <= spriteVisibleReg_32; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1 <= inSpriteHorizontal_32 & inSpriteVertical_32; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_32_REG <= spriteMemories_32_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_33_REG <= spriteMemories_33_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1 <= spriteVisibleReg_33; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1 <= inSpriteHorizontal_33 & inSpriteVertical_33; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_33_REG <= spriteMemories_33_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_34_REG <= spriteMemories_34_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1 <= spriteVisibleReg_34; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1 <= inSpriteHorizontal_34 & inSpriteVertical_34; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_34_REG <= spriteMemories_34_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_35_REG <= spriteMemories_35_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1 <= spriteVisibleReg_35; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1 <= inSpriteHorizontal_35 & inSpriteVertical_35; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_35_REG <= spriteMemories_35_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_36_REG <= spriteMemories_36_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1 <= spriteVisibleReg_36; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1 <= inSpriteHorizontal_36 & inSpriteVertical_36; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_36_REG <= spriteMemories_36_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_37_REG <= spriteMemories_37_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1 <= spriteVisibleReg_37; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1 <= inSpriteHorizontal_37 & inSpriteVertical_37; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_37_REG <= spriteMemories_37_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_38_REG <= spriteMemories_38_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1 <= spriteVisibleReg_38; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1 <= inSpriteHorizontal_38 & inSpriteVertical_38; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_38_REG <= spriteMemories_38_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_39_REG <= spriteMemories_39_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1 <= spriteVisibleReg_39; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1 <= inSpriteHorizontal_39 & inSpriteVertical_39; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_39_REG <= spriteMemories_39_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_40_REG <= spriteMemories_40_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1 <= spriteVisibleReg_40; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1 <= inSpriteHorizontal_40 & inSpriteVertical_40; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_40_REG <= spriteMemories_40_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_41_REG <= spriteMemories_41_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1 <= spriteVisibleReg_41; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1 <= inSpriteHorizontal_41 & inSpriteVertical_41; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_41_REG <= spriteMemories_41_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_42_REG <= spriteMemories_42_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1 <= spriteVisibleReg_42; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1 <= inSpriteHorizontal_42 & inSpriteVertical_42; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_42_REG <= spriteMemories_42_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_43_REG <= spriteMemories_43_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1 <= spriteVisibleReg_43; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1 <= inSpriteHorizontal_43 & inSpriteVertical_43; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_43_REG <= spriteMemories_43_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_44_REG <= spriteMemories_44_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1 <= spriteVisibleReg_44; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1 <= inSpriteHorizontal_44 & inSpriteVertical_44; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_44_REG <= spriteMemories_44_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_45_REG <= spriteMemories_45_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1 <= spriteVisibleReg_45; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1 <= inSpriteHorizontal_45 & inSpriteVertical_45; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_45_REG <= spriteMemories_45_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_46_REG <= spriteMemories_46_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1 <= spriteVisibleReg_46; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1 <= inSpriteHorizontal_46 & inSpriteVertical_46; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_46_REG <= spriteMemories_46_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_47_REG <= spriteMemories_47_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1 <= spriteVisibleReg_47; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1 <= inSpriteHorizontal_47 & inSpriteVertical_47; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_47_REG <= spriteMemories_47_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_48_REG <= spriteMemories_48_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1 <= spriteVisibleReg_48; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1 <= inSpriteHorizontal_48 & inSpriteVertical_48; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_48_REG <= spriteMemories_48_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_49_REG <= spriteMemories_49_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1 <= spriteVisibleReg_49; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1 <= inSpriteHorizontal_49 & inSpriteVertical_49; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_49_REG <= spriteMemories_49_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_50_REG <= spriteMemories_50_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1 <= spriteVisibleReg_50; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1 <= inSpriteHorizontal_50 & inSpriteVertical_50; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_50_REG <= spriteMemories_50_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_51_REG <= spriteMemories_51_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1 <= spriteVisibleReg_51; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1 <= inSpriteHorizontal_51 & inSpriteVertical_51; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_51_REG <= spriteMemories_51_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_52_REG <= spriteMemories_52_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1 <= spriteVisibleReg_52; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1 <= inSpriteHorizontal_52 & inSpriteVertical_52; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_52_REG <= spriteMemories_52_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_53_REG <= spriteMemories_53_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1 <= spriteVisibleReg_53; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1 <= inSpriteHorizontal_53 & inSpriteVertical_53; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_53_REG <= spriteMemories_53_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_54_REG <= spriteMemories_54_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1 <= spriteVisibleReg_54; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1 <= inSpriteHorizontal_54 & inSpriteVertical_54; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_54_REG <= spriteMemories_54_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_55_REG <= spriteMemories_55_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1 <= spriteVisibleReg_55; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1 <= inSpriteHorizontal_55 & inSpriteVertical_55; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_55_REG <= spriteMemories_55_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_56_REG <= spriteMemories_56_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1 <= spriteVisibleReg_56; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1 <= inSpriteHorizontal_56 & inSpriteVertical_56; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_56_REG <= spriteMemories_56_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_57_REG <= spriteMemories_57_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1 <= spriteVisibleReg_57; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1 <= inSpriteHorizontal_57 & inSpriteVertical_57; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_57_REG <= spriteMemories_57_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_58_REG <= spriteMemories_58_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1 <= spriteVisibleReg_58; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1 <= inSpriteHorizontal_58 & inSpriteVertical_58; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_58_REG <= spriteMemories_58_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_59_REG <= spriteMemories_59_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1 <= spriteVisibleReg_59; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1 <= inSpriteHorizontal_59 & inSpriteVertical_59; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_59_REG <= spriteMemories_59_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_60_REG <= spriteMemories_60_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1 <= spriteVisibleReg_60; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1 <= inSpriteHorizontal_60 & inSpriteVertical_60; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_60_REG <= spriteMemories_60_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_61_REG <= spriteMemories_61_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1 <= spriteVisibleReg_61; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1 <= inSpriteHorizontal_61 & inSpriteVertical_61; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_61_REG <= spriteMemories_61_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_62_REG <= spriteMemories_62_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1 <= spriteVisibleReg_62; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1 <= inSpriteHorizontal_62 & inSpriteVertical_62; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_62_REG <= spriteMemories_62_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_63_REG <= spriteMemories_63_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1 <= spriteVisibleReg_63; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1 <= inSpriteHorizontal_63 & inSpriteVertical_63; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_63_REG <= spriteMemories_63_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    pixelColorSprite <= multiHotPriortyReductionTree_io_dataOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 339:33]
    pixelColorSpriteValid <= multiHotPriortyReductionTree_io_selectOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 340:38]
    pixelColourVGA_pipeReg_0 <= pixelColourVGA_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    pixelColourVGA_pipeReg_1 <= pixelColourVGA_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    pixelColourVGA_pipeReg_2 <= CounterXReg < 10'h280 & CounterYReg < 10'h1e0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 97:60]
    io_vgaRed_REG <= {pixelColourVGA[5:4],pixelColourVGA[5:4]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 346:26]
    io_vgaGreen_REG <= {pixelColourVGA[3:2],pixelColourVGA[3:2]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 347:28]
    io_vgaBlue_REG <= {pixelColourVGA[1:0],pixelColourVGA[1:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 348:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ScaleCounterReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  CounterXReg = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  CounterYReg = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  backMemoryRestoreCounter = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  io_Hsync_pipeReg_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_Hsync_pipeReg_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_Hsync_pipeReg_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_Hsync_pipeReg_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_Vsync_pipeReg_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  io_Vsync_pipeReg_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_Vsync_pipeReg_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_Vsync_pipeReg_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  frameClockCount = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXPositionReg_3 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXPositionReg_7 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXPositionReg_8 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXPositionReg_9 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXPositionReg_10 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXPositionReg_11 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXPositionReg_12 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteXPositionReg_13 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  spriteXPositionReg_14 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  spriteXPositionReg_16 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  spriteXPositionReg_17 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  spriteXPositionReg_18 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  spriteXPositionReg_19 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  spriteXPositionReg_20 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  spriteXPositionReg_21 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  spriteXPositionReg_22 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  spriteXPositionReg_23 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  spriteXPositionReg_24 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  spriteXPositionReg_25 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  spriteXPositionReg_26 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  spriteXPositionReg_27 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  spriteXPositionReg_28 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  spriteXPositionReg_29 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  spriteXPositionReg_30 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  spriteXPositionReg_31 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  spriteXPositionReg_32 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  spriteXPositionReg_33 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  spriteXPositionReg_34 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  spriteXPositionReg_35 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  spriteXPositionReg_36 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  spriteXPositionReg_37 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  spriteXPositionReg_38 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  spriteXPositionReg_39 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  spriteXPositionReg_40 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  spriteXPositionReg_41 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  spriteXPositionReg_42 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  spriteXPositionReg_43 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  spriteXPositionReg_44 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  spriteXPositionReg_45 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  spriteXPositionReg_46 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  spriteXPositionReg_47 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  spriteXPositionReg_48 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  spriteXPositionReg_49 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  spriteXPositionReg_50 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  spriteXPositionReg_51 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  spriteXPositionReg_52 = _RAND_58[10:0];
  _RAND_59 = {1{`RANDOM}};
  spriteXPositionReg_53 = _RAND_59[10:0];
  _RAND_60 = {1{`RANDOM}};
  spriteXPositionReg_54 = _RAND_60[10:0];
  _RAND_61 = {1{`RANDOM}};
  spriteXPositionReg_55 = _RAND_61[10:0];
  _RAND_62 = {1{`RANDOM}};
  spriteXPositionReg_56 = _RAND_62[10:0];
  _RAND_63 = {1{`RANDOM}};
  spriteXPositionReg_57 = _RAND_63[10:0];
  _RAND_64 = {1{`RANDOM}};
  spriteXPositionReg_58 = _RAND_64[10:0];
  _RAND_65 = {1{`RANDOM}};
  spriteXPositionReg_59 = _RAND_65[10:0];
  _RAND_66 = {1{`RANDOM}};
  spriteXPositionReg_60 = _RAND_66[10:0];
  _RAND_67 = {1{`RANDOM}};
  spriteXPositionReg_61 = _RAND_67[10:0];
  _RAND_68 = {1{`RANDOM}};
  spriteXPositionReg_62 = _RAND_68[10:0];
  _RAND_69 = {1{`RANDOM}};
  spriteXPositionReg_63 = _RAND_69[10:0];
  _RAND_70 = {1{`RANDOM}};
  spriteYPositionReg_3 = _RAND_70[9:0];
  _RAND_71 = {1{`RANDOM}};
  spriteYPositionReg_7 = _RAND_71[9:0];
  _RAND_72 = {1{`RANDOM}};
  spriteYPositionReg_8 = _RAND_72[9:0];
  _RAND_73 = {1{`RANDOM}};
  spriteYPositionReg_9 = _RAND_73[9:0];
  _RAND_74 = {1{`RANDOM}};
  spriteYPositionReg_10 = _RAND_74[9:0];
  _RAND_75 = {1{`RANDOM}};
  spriteYPositionReg_11 = _RAND_75[9:0];
  _RAND_76 = {1{`RANDOM}};
  spriteYPositionReg_12 = _RAND_76[9:0];
  _RAND_77 = {1{`RANDOM}};
  spriteYPositionReg_13 = _RAND_77[9:0];
  _RAND_78 = {1{`RANDOM}};
  spriteYPositionReg_14 = _RAND_78[9:0];
  _RAND_79 = {1{`RANDOM}};
  spriteYPositionReg_16 = _RAND_79[9:0];
  _RAND_80 = {1{`RANDOM}};
  spriteYPositionReg_17 = _RAND_80[9:0];
  _RAND_81 = {1{`RANDOM}};
  spriteYPositionReg_18 = _RAND_81[9:0];
  _RAND_82 = {1{`RANDOM}};
  spriteYPositionReg_19 = _RAND_82[9:0];
  _RAND_83 = {1{`RANDOM}};
  spriteYPositionReg_20 = _RAND_83[9:0];
  _RAND_84 = {1{`RANDOM}};
  spriteYPositionReg_21 = _RAND_84[9:0];
  _RAND_85 = {1{`RANDOM}};
  spriteYPositionReg_22 = _RAND_85[9:0];
  _RAND_86 = {1{`RANDOM}};
  spriteYPositionReg_23 = _RAND_86[9:0];
  _RAND_87 = {1{`RANDOM}};
  spriteYPositionReg_24 = _RAND_87[9:0];
  _RAND_88 = {1{`RANDOM}};
  spriteYPositionReg_25 = _RAND_88[9:0];
  _RAND_89 = {1{`RANDOM}};
  spriteYPositionReg_26 = _RAND_89[9:0];
  _RAND_90 = {1{`RANDOM}};
  spriteYPositionReg_27 = _RAND_90[9:0];
  _RAND_91 = {1{`RANDOM}};
  spriteYPositionReg_28 = _RAND_91[9:0];
  _RAND_92 = {1{`RANDOM}};
  spriteYPositionReg_29 = _RAND_92[9:0];
  _RAND_93 = {1{`RANDOM}};
  spriteYPositionReg_30 = _RAND_93[9:0];
  _RAND_94 = {1{`RANDOM}};
  spriteYPositionReg_31 = _RAND_94[9:0];
  _RAND_95 = {1{`RANDOM}};
  spriteYPositionReg_32 = _RAND_95[9:0];
  _RAND_96 = {1{`RANDOM}};
  spriteYPositionReg_33 = _RAND_96[9:0];
  _RAND_97 = {1{`RANDOM}};
  spriteYPositionReg_34 = _RAND_97[9:0];
  _RAND_98 = {1{`RANDOM}};
  spriteYPositionReg_35 = _RAND_98[9:0];
  _RAND_99 = {1{`RANDOM}};
  spriteYPositionReg_36 = _RAND_99[9:0];
  _RAND_100 = {1{`RANDOM}};
  spriteYPositionReg_37 = _RAND_100[9:0];
  _RAND_101 = {1{`RANDOM}};
  spriteYPositionReg_38 = _RAND_101[9:0];
  _RAND_102 = {1{`RANDOM}};
  spriteYPositionReg_39 = _RAND_102[9:0];
  _RAND_103 = {1{`RANDOM}};
  spriteYPositionReg_40 = _RAND_103[9:0];
  _RAND_104 = {1{`RANDOM}};
  spriteYPositionReg_41 = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  spriteYPositionReg_42 = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  spriteYPositionReg_43 = _RAND_106[9:0];
  _RAND_107 = {1{`RANDOM}};
  spriteYPositionReg_44 = _RAND_107[9:0];
  _RAND_108 = {1{`RANDOM}};
  spriteYPositionReg_45 = _RAND_108[9:0];
  _RAND_109 = {1{`RANDOM}};
  spriteYPositionReg_46 = _RAND_109[9:0];
  _RAND_110 = {1{`RANDOM}};
  spriteYPositionReg_47 = _RAND_110[9:0];
  _RAND_111 = {1{`RANDOM}};
  spriteYPositionReg_48 = _RAND_111[9:0];
  _RAND_112 = {1{`RANDOM}};
  spriteYPositionReg_49 = _RAND_112[9:0];
  _RAND_113 = {1{`RANDOM}};
  spriteYPositionReg_50 = _RAND_113[9:0];
  _RAND_114 = {1{`RANDOM}};
  spriteYPositionReg_51 = _RAND_114[9:0];
  _RAND_115 = {1{`RANDOM}};
  spriteYPositionReg_52 = _RAND_115[9:0];
  _RAND_116 = {1{`RANDOM}};
  spriteYPositionReg_53 = _RAND_116[9:0];
  _RAND_117 = {1{`RANDOM}};
  spriteYPositionReg_54 = _RAND_117[9:0];
  _RAND_118 = {1{`RANDOM}};
  spriteYPositionReg_55 = _RAND_118[9:0];
  _RAND_119 = {1{`RANDOM}};
  spriteYPositionReg_56 = _RAND_119[9:0];
  _RAND_120 = {1{`RANDOM}};
  spriteYPositionReg_57 = _RAND_120[9:0];
  _RAND_121 = {1{`RANDOM}};
  spriteYPositionReg_58 = _RAND_121[9:0];
  _RAND_122 = {1{`RANDOM}};
  spriteYPositionReg_59 = _RAND_122[9:0];
  _RAND_123 = {1{`RANDOM}};
  spriteYPositionReg_60 = _RAND_123[9:0];
  _RAND_124 = {1{`RANDOM}};
  spriteYPositionReg_61 = _RAND_124[9:0];
  _RAND_125 = {1{`RANDOM}};
  spriteYPositionReg_62 = _RAND_125[9:0];
  _RAND_126 = {1{`RANDOM}};
  spriteYPositionReg_63 = _RAND_126[9:0];
  _RAND_127 = {1{`RANDOM}};
  spriteVisibleReg_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  spriteVisibleReg_1 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  spriteVisibleReg_2 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  spriteVisibleReg_3 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  spriteVisibleReg_4 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  spriteVisibleReg_5 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  spriteVisibleReg_6 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  spriteVisibleReg_7 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  spriteVisibleReg_8 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  spriteVisibleReg_9 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  spriteVisibleReg_10 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  spriteVisibleReg_11 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  spriteVisibleReg_12 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  spriteVisibleReg_13 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  spriteVisibleReg_14 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  spriteVisibleReg_15 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  spriteVisibleReg_16 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  spriteVisibleReg_17 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  spriteVisibleReg_18 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  spriteVisibleReg_19 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  spriteVisibleReg_20 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  spriteVisibleReg_21 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  spriteVisibleReg_22 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  spriteVisibleReg_23 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  spriteVisibleReg_24 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  spriteVisibleReg_25 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  spriteVisibleReg_26 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  spriteVisibleReg_27 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  spriteVisibleReg_28 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  spriteVisibleReg_29 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  spriteVisibleReg_30 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  spriteVisibleReg_31 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  spriteVisibleReg_32 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  spriteVisibleReg_33 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  spriteVisibleReg_34 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  spriteVisibleReg_35 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  spriteVisibleReg_36 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  spriteVisibleReg_37 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  spriteVisibleReg_38 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  spriteVisibleReg_39 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  spriteVisibleReg_40 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  spriteVisibleReg_41 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  spriteVisibleReg_42 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  spriteVisibleReg_43 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  spriteVisibleReg_44 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  spriteVisibleReg_45 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  spriteVisibleReg_46 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  spriteVisibleReg_47 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  spriteVisibleReg_48 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  spriteVisibleReg_49 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  spriteVisibleReg_50 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  spriteVisibleReg_51 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  spriteVisibleReg_52 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  spriteVisibleReg_53 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  spriteVisibleReg_54 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  spriteVisibleReg_55 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  spriteVisibleReg_56 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  spriteVisibleReg_57 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  spriteVisibleReg_58 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  spriteVisibleReg_59 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  spriteVisibleReg_60 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  spriteVisibleReg_61 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  spriteVisibleReg_62 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  spriteVisibleReg_63 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_16 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_17 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_18 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_19 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_20 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_21 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_22 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_23 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_24 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_25 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_26 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_27 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_28 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_29 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_30 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_31 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_32 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_33 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_34 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_35 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_36 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_37 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_38 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_39 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_40 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_41 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_42 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_43 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_44 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_45 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_58 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_59 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  spriteScaleUpHorizontalReg_60 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_16 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_17 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_18 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_19 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_20 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_21 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_22 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_23 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_24 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_25 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_26 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_27 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_28 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_29 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_30 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_31 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_32 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_33 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_34 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_35 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_36 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_37 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_38 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_39 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_40 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_41 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_42 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_43 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_44 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_45 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_58 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_59 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  spriteScaleUpVerticalReg_60 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  viewBoxXReg = _RAND_257[9:0];
  _RAND_258 = {1{`RANDOM}};
  viewBoxYReg = _RAND_258[8:0];
  _RAND_259 = {1{`RANDOM}};
  missingFrameErrorReg = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  viewBoxOutOfRangeErrorReg = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  newFrameStikyReg = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  REG = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  backTileMemoryDataRead_0_REG = _RAND_263[6:0];
  _RAND_264 = {1{`RANDOM}};
  backTileMemoryDataRead_1_REG = _RAND_264[6:0];
  _RAND_265 = {1{`RANDOM}};
  backTileMemoryDataRead_2_REG = _RAND_265[6:0];
  _RAND_266 = {1{`RANDOM}};
  backTileMemoryDataRead_3_REG = _RAND_266[6:0];
  _RAND_267 = {1{`RANDOM}};
  backTileMemoryDataRead_4_REG = _RAND_267[6:0];
  _RAND_268 = {1{`RANDOM}};
  backTileMemoryDataRead_5_REG = _RAND_268[6:0];
  _RAND_269 = {1{`RANDOM}};
  backTileMemoryDataRead_6_REG = _RAND_269[6:0];
  _RAND_270 = {1{`RANDOM}};
  backTileMemoryDataRead_7_REG = _RAND_270[6:0];
  _RAND_271 = {1{`RANDOM}};
  backTileMemoryDataRead_8_REG = _RAND_271[6:0];
  _RAND_272 = {1{`RANDOM}};
  backTileMemoryDataRead_9_REG = _RAND_272[6:0];
  _RAND_273 = {1{`RANDOM}};
  backTileMemoryDataRead_10_REG = _RAND_273[6:0];
  _RAND_274 = {1{`RANDOM}};
  backTileMemoryDataRead_11_REG = _RAND_274[6:0];
  _RAND_275 = {1{`RANDOM}};
  backTileMemoryDataRead_12_REG = _RAND_275[6:0];
  _RAND_276 = {1{`RANDOM}};
  backTileMemoryDataRead_13_REG = _RAND_276[6:0];
  _RAND_277 = {1{`RANDOM}};
  backTileMemoryDataRead_14_REG = _RAND_277[6:0];
  _RAND_278 = {1{`RANDOM}};
  backTileMemoryDataRead_15_REG = _RAND_278[6:0];
  _RAND_279 = {1{`RANDOM}};
  backTileMemoryDataRead_16_REG = _RAND_279[6:0];
  _RAND_280 = {1{`RANDOM}};
  backTileMemoryDataRead_17_REG = _RAND_280[6:0];
  _RAND_281 = {1{`RANDOM}};
  backTileMemoryDataRead_18_REG = _RAND_281[6:0];
  _RAND_282 = {1{`RANDOM}};
  backTileMemoryDataRead_19_REG = _RAND_282[6:0];
  _RAND_283 = {1{`RANDOM}};
  backTileMemoryDataRead_20_REG = _RAND_283[6:0];
  _RAND_284 = {1{`RANDOM}};
  backTileMemoryDataRead_21_REG = _RAND_284[6:0];
  _RAND_285 = {1{`RANDOM}};
  backTileMemoryDataRead_22_REG = _RAND_285[6:0];
  _RAND_286 = {1{`RANDOM}};
  backTileMemoryDataRead_23_REG = _RAND_286[6:0];
  _RAND_287 = {1{`RANDOM}};
  backTileMemoryDataRead_24_REG = _RAND_287[6:0];
  _RAND_288 = {1{`RANDOM}};
  backTileMemoryDataRead_25_REG = _RAND_288[6:0];
  _RAND_289 = {1{`RANDOM}};
  backTileMemoryDataRead_26_REG = _RAND_289[6:0];
  _RAND_290 = {1{`RANDOM}};
  backTileMemoryDataRead_27_REG = _RAND_290[6:0];
  _RAND_291 = {1{`RANDOM}};
  backTileMemoryDataRead_28_REG = _RAND_291[6:0];
  _RAND_292 = {1{`RANDOM}};
  backTileMemoryDataRead_29_REG = _RAND_292[6:0];
  _RAND_293 = {1{`RANDOM}};
  backTileMemoryDataRead_30_REG = _RAND_293[6:0];
  _RAND_294 = {1{`RANDOM}};
  backTileMemoryDataRead_31_REG = _RAND_294[6:0];
  _RAND_295 = {1{`RANDOM}};
  backTileMemoryDataRead_32_REG = _RAND_295[6:0];
  _RAND_296 = {1{`RANDOM}};
  backTileMemoryDataRead_33_REG = _RAND_296[6:0];
  _RAND_297 = {1{`RANDOM}};
  backTileMemoryDataRead_34_REG = _RAND_297[6:0];
  _RAND_298 = {1{`RANDOM}};
  backTileMemoryDataRead_35_REG = _RAND_298[6:0];
  _RAND_299 = {1{`RANDOM}};
  backTileMemoryDataRead_36_REG = _RAND_299[6:0];
  _RAND_300 = {1{`RANDOM}};
  backTileMemoryDataRead_37_REG = _RAND_300[6:0];
  _RAND_301 = {1{`RANDOM}};
  backTileMemoryDataRead_38_REG = _RAND_301[6:0];
  _RAND_302 = {1{`RANDOM}};
  backTileMemoryDataRead_39_REG = _RAND_302[6:0];
  _RAND_303 = {1{`RANDOM}};
  backTileMemoryDataRead_40_REG = _RAND_303[6:0];
  _RAND_304 = {1{`RANDOM}};
  backTileMemoryDataRead_41_REG = _RAND_304[6:0];
  _RAND_305 = {1{`RANDOM}};
  backTileMemoryDataRead_42_REG = _RAND_305[6:0];
  _RAND_306 = {1{`RANDOM}};
  backTileMemoryDataRead_43_REG = _RAND_306[6:0];
  _RAND_307 = {1{`RANDOM}};
  backTileMemoryDataRead_44_REG = _RAND_307[6:0];
  _RAND_308 = {1{`RANDOM}};
  backTileMemoryDataRead_45_REG = _RAND_308[6:0];
  _RAND_309 = {1{`RANDOM}};
  backTileMemoryDataRead_46_REG = _RAND_309[6:0];
  _RAND_310 = {1{`RANDOM}};
  backTileMemoryDataRead_47_REG = _RAND_310[6:0];
  _RAND_311 = {1{`RANDOM}};
  backTileMemoryDataRead_48_REG = _RAND_311[6:0];
  _RAND_312 = {1{`RANDOM}};
  backTileMemoryDataRead_49_REG = _RAND_312[6:0];
  _RAND_313 = {1{`RANDOM}};
  backTileMemoryDataRead_50_REG = _RAND_313[6:0];
  _RAND_314 = {1{`RANDOM}};
  backTileMemoryDataRead_51_REG = _RAND_314[6:0];
  _RAND_315 = {1{`RANDOM}};
  backTileMemoryDataRead_52_REG = _RAND_315[6:0];
  _RAND_316 = {1{`RANDOM}};
  backTileMemoryDataRead_53_REG = _RAND_316[6:0];
  _RAND_317 = {1{`RANDOM}};
  backTileMemoryDataRead_54_REG = _RAND_317[6:0];
  _RAND_318 = {1{`RANDOM}};
  backTileMemoryDataRead_55_REG = _RAND_318[6:0];
  _RAND_319 = {1{`RANDOM}};
  backTileMemoryDataRead_56_REG = _RAND_319[6:0];
  _RAND_320 = {1{`RANDOM}};
  backTileMemoryDataRead_57_REG = _RAND_320[6:0];
  _RAND_321 = {1{`RANDOM}};
  backTileMemoryDataRead_58_REG = _RAND_321[6:0];
  _RAND_322 = {1{`RANDOM}};
  backTileMemoryDataRead_59_REG = _RAND_322[6:0];
  _RAND_323 = {1{`RANDOM}};
  backTileMemoryDataRead_60_REG = _RAND_323[6:0];
  _RAND_324 = {1{`RANDOM}};
  backTileMemoryDataRead_61_REG = _RAND_324[6:0];
  _RAND_325 = {1{`RANDOM}};
  backTileMemoryDataRead_62_REG = _RAND_325[6:0];
  _RAND_326 = {1{`RANDOM}};
  backTileMemoryDataRead_63_REG = _RAND_326[6:0];
  _RAND_327 = {1{`RANDOM}};
  backMemoryCopyCounter = _RAND_327[11:0];
  _RAND_328 = {1{`RANDOM}};
  copyEnabledReg = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  backBufferShadowMemory_io_address_REG = _RAND_329[10:0];
  _RAND_330 = {1{`RANDOM}};
  backBufferShadowMemory_io_writeEnable_REG = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  backBufferMemory_io_address_REG = _RAND_331[10:0];
  _RAND_332 = {1{`RANDOM}};
  fullBackgroundColor_REG = _RAND_332[5:0];
  _RAND_333 = {1{`RANDOM}};
  pixelColorBack = _RAND_333[5:0];
  _RAND_334 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_0_REG = _RAND_334[5:0];
  _RAND_335 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_REG = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_1_REG = _RAND_340[5:0];
  _RAND_341 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_REG = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_2_REG = _RAND_346[5:0];
  _RAND_347 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_REG = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_3_REG = _RAND_352[5:0];
  _RAND_353 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_REG = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_4_REG = _RAND_358[5:0];
  _RAND_359 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_REG = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_5_REG = _RAND_364[5:0];
  _RAND_365 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_REG = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_6_REG = _RAND_370[5:0];
  _RAND_371 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_REG = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_7_REG = _RAND_376[5:0];
  _RAND_377 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_REG = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_8_REG = _RAND_382[5:0];
  _RAND_383 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_REG = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_9_REG = _RAND_388[5:0];
  _RAND_389 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_REG = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_10_REG = _RAND_394[5:0];
  _RAND_395 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_REG = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_11_REG = _RAND_400[5:0];
  _RAND_401 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_REG = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_12_REG = _RAND_406[5:0];
  _RAND_407 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_REG = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_13_REG = _RAND_412[5:0];
  _RAND_413 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_REG = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_14_REG = _RAND_418[5:0];
  _RAND_419 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_REG = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_15_REG = _RAND_424[5:0];
  _RAND_425 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_REG = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_16_REG = _RAND_430[5:0];
  _RAND_431 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_REG = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_17_REG = _RAND_436[5:0];
  _RAND_437 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_REG = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_18_REG = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_REG = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_19_REG = _RAND_448[5:0];
  _RAND_449 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_REG = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_20_REG = _RAND_454[5:0];
  _RAND_455 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_REG = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_21_REG = _RAND_460[5:0];
  _RAND_461 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_REG = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_22_REG = _RAND_466[5:0];
  _RAND_467 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_REG = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_23_REG = _RAND_472[5:0];
  _RAND_473 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_REG = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_24_REG = _RAND_478[5:0];
  _RAND_479 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_REG = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_25_REG = _RAND_484[5:0];
  _RAND_485 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_REG = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_26_REG = _RAND_490[5:0];
  _RAND_491 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_REG = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_27_REG = _RAND_496[5:0];
  _RAND_497 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_REG = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_28_REG = _RAND_502[5:0];
  _RAND_503 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_REG = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_29_REG = _RAND_508[5:0];
  _RAND_509 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_REG = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_30_REG = _RAND_514[5:0];
  _RAND_515 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_REG = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_31_REG = _RAND_520[5:0];
  _RAND_521 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_REG = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_32_REG = _RAND_526[5:0];
  _RAND_527 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__0 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg__1 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_0 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_pipeReg_1_1 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_32_REG = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_33_REG = _RAND_532[5:0];
  _RAND_533 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__0 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg__1 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_0 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_pipeReg_1_1 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_33_REG = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_34_REG = _RAND_538[5:0];
  _RAND_539 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__0 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg__1 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_0 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_pipeReg_1_1 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_34_REG = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_35_REG = _RAND_544[5:0];
  _RAND_545 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__0 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg__1 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_0 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_pipeReg_1_1 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_35_REG = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_36_REG = _RAND_550[5:0];
  _RAND_551 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__0 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg__1 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_0 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_pipeReg_1_1 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_36_REG = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_37_REG = _RAND_556[5:0];
  _RAND_557 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__0 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg__1 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_0 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_pipeReg_1_1 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_37_REG = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_38_REG = _RAND_562[5:0];
  _RAND_563 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__0 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg__1 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_0 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_pipeReg_1_1 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_38_REG = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_39_REG = _RAND_568[5:0];
  _RAND_569 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__0 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg__1 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_0 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_pipeReg_1_1 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_39_REG = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_40_REG = _RAND_574[5:0];
  _RAND_575 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__0 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg__1 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_0 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_pipeReg_1_1 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_40_REG = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_41_REG = _RAND_580[5:0];
  _RAND_581 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__0 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg__1 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_0 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_pipeReg_1_1 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_41_REG = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_42_REG = _RAND_586[5:0];
  _RAND_587 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__0 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg__1 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_0 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_pipeReg_1_1 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_42_REG = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_43_REG = _RAND_592[5:0];
  _RAND_593 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__0 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg__1 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_0 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_pipeReg_1_1 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_43_REG = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_44_REG = _RAND_598[5:0];
  _RAND_599 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__0 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg__1 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_0 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_pipeReg_1_1 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_44_REG = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_45_REG = _RAND_604[5:0];
  _RAND_605 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__0 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg__1 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_0 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_pipeReg_1_1 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_45_REG = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_46_REG = _RAND_610[5:0];
  _RAND_611 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__0 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg__1 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_0 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_pipeReg_1_1 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_46_REG = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_47_REG = _RAND_616[5:0];
  _RAND_617 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__0 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg__1 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_0 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_pipeReg_1_1 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_47_REG = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_48_REG = _RAND_622[5:0];
  _RAND_623 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__0 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg__1 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_0 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_pipeReg_1_1 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_48_REG = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_49_REG = _RAND_628[5:0];
  _RAND_629 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__0 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg__1 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_0 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_pipeReg_1_1 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_49_REG = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_50_REG = _RAND_634[5:0];
  _RAND_635 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__0 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg__1 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_0 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_pipeReg_1_1 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_50_REG = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_51_REG = _RAND_640[5:0];
  _RAND_641 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__0 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg__1 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_0 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_pipeReg_1_1 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_51_REG = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_52_REG = _RAND_646[5:0];
  _RAND_647 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__0 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg__1 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_0 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_pipeReg_1_1 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_52_REG = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_53_REG = _RAND_652[5:0];
  _RAND_653 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__0 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg__1 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_0 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_pipeReg_1_1 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_53_REG = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_54_REG = _RAND_658[5:0];
  _RAND_659 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__0 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg__1 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_0 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_pipeReg_1_1 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_54_REG = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_55_REG = _RAND_664[5:0];
  _RAND_665 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__0 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg__1 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_0 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_pipeReg_1_1 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_55_REG = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_56_REG = _RAND_670[5:0];
  _RAND_671 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__0 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg__1 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_0 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_pipeReg_1_1 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_56_REG = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_57_REG = _RAND_676[5:0];
  _RAND_677 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__0 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg__1 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_0 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_pipeReg_1_1 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_57_REG = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_58_REG = _RAND_682[5:0];
  _RAND_683 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__0 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg__1 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_0 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_pipeReg_1_1 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_58_REG = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_59_REG = _RAND_688[5:0];
  _RAND_689 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__0 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg__1 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_0 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_pipeReg_1_1 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_59_REG = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_60_REG = _RAND_694[5:0];
  _RAND_695 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__0 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg__1 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_0 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_pipeReg_1_1 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_60_REG = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_61_REG = _RAND_700[5:0];
  _RAND_701 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__0 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg__1 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_0 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_pipeReg_1_1 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_61_REG = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_62_REG = _RAND_706[5:0];
  _RAND_707 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__0 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg__1 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_0 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_pipeReg_1_1 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_62_REG = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_63_REG = _RAND_712[5:0];
  _RAND_713 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__0 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg__1 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_0 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_pipeReg_1_1 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_63_REG = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  pixelColorSprite = _RAND_718[5:0];
  _RAND_719 = {1{`RANDOM}};
  pixelColorSpriteValid = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_0 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_1 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_2 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  io_vgaRed_REG = _RAND_723[3:0];
  _RAND_724 = {1{`RANDOM}};
  io_vgaGreen_REG = _RAND_724[3:0];
  _RAND_725 = {1{`RANDOM}};
  io_vgaBlue_REG = _RAND_725[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Memory_131(
  input         clock,
  input  [7:0]  io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [27:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [7:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(8), .DATA_WIDTH(28), .LOAD_FILE("memory_init/tune_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 28'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_132(
  input         clock,
  input  [7:0]  io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [27:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [7:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(8), .DATA_WIDTH(28), .LOAD_FILE("memory_init/tune_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 28'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module SoundEngine(
  input   clock,
  input   reset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  tuneMemories_0_clock; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [7:0] tuneMemories_0_io_address; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [27:0] tuneMemories_0_io_dataRead; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire  tuneMemories_1_clock; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [7:0] tuneMemories_1_io_address; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [27:0] tuneMemories_1_io_dataRead; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  reg [11:0] durationCountReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
  reg [11:0] durationCountReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
  reg [11:0] currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
  reg [11:0] currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
  reg [7:0] nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
  reg [7:0] nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
  reg [1:0] stateReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
  reg [1:0] stateReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
  reg  newNoteLoadReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
  reg  newNoteLoadReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
  wire  durationCountRegDone_0 = durationCountReg_0 == 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 89:54]
  wire  _T_8 = tuneMemories_0_io_dataRead[27:16] != 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 111:60]
  wire [1:0] _GEN_4 = tuneMemories_0_io_dataRead[27:16] != 12'h0 ? 2'h3 : stateReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 112:23 62:25]
  wire [11:0] _GEN_6 = tuneMemories_0_io_dataRead[27:16] != 12'h0 ? tuneMemories_0_io_dataRead[27:16] :
    currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 114:30 58:32]
  wire  _T_13 = durationCountRegDone_0 & ~newNoteLoadReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:44]
  wire [7:0] _nextIndexReg_0_T_1 = nextIndexReg_0 + 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 126:46]
  wire [11:0] _GEN_10 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? tuneMemories_0_io_dataRead[27:16] :
    currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 124:30 58:32]
  wire [7:0] _GEN_12 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? _nextIndexReg_0_T_1 : nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 126:27 59:29]
  wire [7:0] _GEN_14 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? 8'h0 : _GEN_12; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 120:27]
  wire [11:0] _GEN_16 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? currDurationReg_0 : _GEN_10; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 58:32]
  wire  _GEN_17 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? 1'h0 : _T_13; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 97:23]
  wire [7:0] _GEN_22 = 2'h3 == stateReg_0 ? _GEN_14 : nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 59:29]
  wire [11:0] _GEN_24 = 2'h3 == stateReg_0 ? _GEN_16 : currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 58:32]
  wire  _GEN_25 = 2'h3 == stateReg_0 & _GEN_17; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 97:23]
  wire  durationCountRegDone_1 = durationCountReg_1 == 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 89:54]
  wire  _T_25 = tuneMemories_1_io_dataRead[27:16] != 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 111:60]
  wire [1:0] _GEN_52 = tuneMemories_1_io_dataRead[27:16] != 12'h0 ? 2'h3 : stateReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 112:23 62:25]
  wire [11:0] _GEN_54 = tuneMemories_1_io_dataRead[27:16] != 12'h0 ? tuneMemories_1_io_dataRead[27:16] :
    currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 114:30 58:32]
  wire  _T_30 = durationCountRegDone_1 & ~newNoteLoadReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:44]
  wire [7:0] _nextIndexReg_1_T_1 = nextIndexReg_1 + 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 126:46]
  wire [11:0] _GEN_58 = durationCountRegDone_1 & ~newNoteLoadReg_1 ? tuneMemories_1_io_dataRead[27:16] :
    currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 124:30 58:32]
  wire [7:0] _GEN_60 = durationCountRegDone_1 & ~newNoteLoadReg_1 ? _nextIndexReg_1_T_1 : nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 126:27 59:29]
  wire [7:0] _GEN_62 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? 8'h0 : _GEN_60; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 120:27]
  wire [11:0] _GEN_64 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? currDurationReg_1 : _GEN_58; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 58:32]
  wire  _GEN_65 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? 1'h0 : _T_30; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 97:23]
  wire [7:0] _GEN_70 = 2'h3 == stateReg_1 ? _GEN_62 : nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 59:29]
  wire [11:0] _GEN_72 = 2'h3 == stateReg_1 ? _GEN_64 : currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 58:32]
  wire  _GEN_73 = 2'h3 == stateReg_1 & _GEN_65; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 97:23]
  Memory_131 tuneMemories_0 ( // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
    .clock(tuneMemories_0_clock),
    .io_address(tuneMemories_0_io_address),
    .io_dataRead(tuneMemories_0_io_dataRead)
  );
  Memory_132 tuneMemories_1 ( // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
    .clock(tuneMemories_1_clock),
    .io_address(tuneMemories_1_io_address),
    .io_dataRead(tuneMemories_1_io_dataRead)
  );
  assign tuneMemories_0_clock = clock;
  assign tuneMemories_0_io_address = nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 72:32]
  assign tuneMemories_1_clock = clock;
  assign tuneMemories_1_io_address = nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 72:32]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
      durationCountReg_0 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
    end else if (newNoteLoadReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 84:35]
      durationCountReg_0 <= currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 85:27]
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
      durationCountReg_1 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
    end else if (newNoteLoadReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 84:35]
      durationCountReg_1 <= currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 85:27]
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
      currDurationReg_0 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
    end else if (!(2'h0 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h1 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
          currDurationReg_0 <= _GEN_6;
        end else begin
          currDurationReg_0 <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
      currDurationReg_1 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
    end else if (!(2'h0 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h1 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
          currDurationReg_1 <= _GEN_54;
        end else begin
          currDurationReg_1 <= _GEN_72;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
      nextIndexReg_0 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 102:25]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 107:25]
    end else if (!(2'h2 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= _GEN_22;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
      nextIndexReg_1 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 102:25]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 107:25]
    end else if (!(2'h2 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= _GEN_70;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
      stateReg_0 <= 2'h0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= 2'h1; // @[\\src\\main\\scala\\SoundEngine.scala 103:21]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= 2'h2; // @[\\src\\main\\scala\\SoundEngine.scala 108:21]
    end else if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= _GEN_4;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
      stateReg_1 <= 2'h0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= 2'h1; // @[\\src\\main\\scala\\SoundEngine.scala 103:21]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= 2'h2; // @[\\src\\main\\scala\\SoundEngine.scala 108:21]
    end else if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= _GEN_52;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= _T_8;
    end else begin
      newNoteLoadReg_0 <= _GEN_25;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= _T_25;
    end else begin
      newNoteLoadReg_1 <= _GEN_73;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  durationCountReg_0 = _RAND_0[11:0];
  _RAND_1 = {1{`RANDOM}};
  durationCountReg_1 = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  currDurationReg_0 = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  currDurationReg_1 = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  nextIndexReg_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  nextIndexReg_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  stateReg_0 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  stateReg_1 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  newNoteLoadReg_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  newNoteLoadReg_1 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Difficulty(
  input         clock,
  input         reset,
  input  [1:0]  io_level, // @[\\src\\main\\scala\\Difficulty.scala 5:14]
  output [26:0] io_speed, // @[\\src\\main\\scala\\Difficulty.scala 5:14]
  input         io_resetSpeed // @[\\src\\main\\scala\\Difficulty.scala 5:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [26:0] speedCnt; // @[\\src\\main\\scala\\Difficulty.scala 13:25]
  reg [26:0] frameDivider; // @[\\src\\main\\scala\\Difficulty.scala 16:29]
  wire  tick = frameDivider == 27'h196e6a; // @[\\src\\main\\scala\\Difficulty.scala 23:21]
  wire [26:0] _frameDivider_T_1 = frameDivider + 27'h1; // @[\\src\\main\\scala\\Difficulty.scala 27:34]
  wire [26:0] _speedCnt_T_1 = speedCnt + 27'h1; // @[\\src\\main\\scala\\Difficulty.scala 34:26]
  wire [22:0] timeInSeconds = speedCnt[26:4]; // @[\\src\\main\\scala\\Difficulty.scala 39:32]
  wire [19:0] scaledTime = timeInSeconds[22:3]; // @[\\src\\main\\scala\\Difficulty.scala 40:34]
  wire  _speedFactor_T = 2'h1 == io_level; // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [1:0] _speedFactor_T_1 = 2'h1 == io_level ? $signed(2'sh1) : $signed(2'sh0); // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire  _speedFactor_T_2 = 2'h2 == io_level; // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [1:0] _speedFactor_T_3 = 2'h2 == io_level ? $signed(2'sh1) : $signed(_speedFactor_T_1); // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire  _speedFactor_T_4 = 2'h3 == io_level; // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [2:0] speedFactor = 2'h3 == io_level ? $signed(3'sh2) : $signed({{1{_speedFactor_T_3[1]}},_speedFactor_T_3}); // @[\\src\\main\\scala\\Difficulty.scala 42:45]
  wire [39:0] _rawSpeed_T = scaledTime * scaledTime; // @[\\src\\main\\scala\\Difficulty.scala 48:37]
  wire [42:0] _rawSpeed_T_1 = $signed(_rawSpeed_T) * $signed(speedFactor); // @[\\src\\main\\scala\\Difficulty.scala 48:44]
  wire [42:0] rawSpeed = 43'sh2 + $signed(_rawSpeed_T_1); // @[\\src\\main\\scala\\Difficulty.scala 48:22]
  wire [4:0] _speedCap_T_1 = _speedFactor_T ? $signed(5'shc) : $signed(5'sha); // @[\\src\\main\\scala\\Difficulty.scala 50:43]
  wire [5:0] _speedCap_T_3 = _speedFactor_T_2 ? $signed(6'sh10) : $signed({{1{_speedCap_T_1[4]}},_speedCap_T_1}); // @[\\src\\main\\scala\\Difficulty.scala 50:43]
  wire [5:0] speedCap = _speedFactor_T_4 ? $signed(6'sh16) : $signed(_speedCap_T_3); // @[\\src\\main\\scala\\Difficulty.scala 50:43]
  wire [42:0] _GEN_4 = {{37{speedCap[5]}},speedCap}; // @[\\src\\main\\scala\\Difficulty.scala 55:28]
  wire [42:0] _io_speed_T_1 = $signed(rawSpeed) > $signed(_GEN_4) ? $signed({{37{speedCap[5]}},speedCap}) : $signed(
    rawSpeed); // @[\\src\\main\\scala\\Difficulty.scala 55:18]
  assign io_speed = _io_speed_T_1[26:0]; // @[\\src\\main\\scala\\Difficulty.scala 55:12]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\Difficulty.scala 13:25]
      speedCnt <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 13:25]
    end else if (io_resetSpeed) begin // @[\\src\\main\\scala\\Difficulty.scala 31:23]
      speedCnt <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 32:14]
    end else if (tick) begin // @[\\src\\main\\scala\\Difficulty.scala 33:20]
      speedCnt <= _speedCnt_T_1; // @[\\src\\main\\scala\\Difficulty.scala 34:14]
    end
    if (reset) begin // @[\\src\\main\\scala\\Difficulty.scala 16:29]
      frameDivider <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 16:29]
    end else if (tick) begin // @[\\src\\main\\scala\\Difficulty.scala 23:37]
      frameDivider <= 27'h0; // @[\\src\\main\\scala\\Difficulty.scala 24:18]
    end else begin
      frameDivider <= _frameDivider_T_1; // @[\\src\\main\\scala\\Difficulty.scala 27:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  speedCnt = _RAND_0[26:0];
  _RAND_1 = {1{`RANDOM}};
  frameDivider = _RAND_1[26:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LFSR(
  input        clock,
  input        reset,
  output [9:0] io_out_0, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_1, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_2, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_3, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_4, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_5, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_6, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_7, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_8, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_9, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_10, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_11, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_12, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_13, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_14, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_15, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_16, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_17, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_18, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_19, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_20, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_21, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_22, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_23, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_24, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_25, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_26, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_27, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_28, // @[\\src\\main\\scala\\LFSR.scala 5:14]
  output [9:0] io_out_29 // @[\\src\\main\\scala\\LFSR.scala 5:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] reg_; // @[\\src\\main\\scala\\LFSR.scala 10:20]
  wire  feedback = reg_[63] ^ reg_[62] ^ reg_[60] ^ reg_[59]; // @[\\src\\main\\scala\\LFSR.scala 13:46]
  wire [63:0] _reg_T_1 = {reg_[62:0],feedback}; // @[\\src\\main\\scala\\LFSR.scala 16:13]
  wire [8:0] current_output = reg_[17:9]; // @[\\src\\main\\scala\\LFSR.scala 19:27]
  reg [9:0] history_0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_1; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_2; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_3; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_4; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_5; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_6; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_7; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_8; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_9; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_10; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_11; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_12; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_13; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_14; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_15; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_16; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_17; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_18; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_19; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_20; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_21; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_22; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_23; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_24; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_25; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_26; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_27; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_28; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  reg [9:0] history_29; // @[\\src\\main\\scala\\LFSR.scala 22:24]
  assign io_out_0 = history_0; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_1 = history_1; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_2 = history_2; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_3 = history_3; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_4 = history_4; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_5 = history_5; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_6 = history_6; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_7 = history_7; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_8 = history_8; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_9 = history_9; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_10 = history_10; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_11 = history_11; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_12 = history_12; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_13 = history_13; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_14 = history_14; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_15 = history_15; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_16 = history_16; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_17 = history_17; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_18 = history_18; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_19 = history_19; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_20 = history_20; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_21 = history_21; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_22 = history_22; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_23 = history_23; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_24 = history_24; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_25 = history_25; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_26 = history_26; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_27 = history_27; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_28 = history_28; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  assign io_out_29 = history_29; // @[\\src\\main\\scala\\LFSR.scala 30:10]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 10:20]
      reg_ <= 64'h123456789abcdef; // @[\\src\\main\\scala\\LFSR.scala 10:20]
    end else begin
      reg_ <= _reg_T_1; // @[\\src\\main\\scala\\LFSR.scala 16:7]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_0 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_0 <= history_1; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_1 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_1 <= history_2; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_2 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_2 <= history_3; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_3 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_3 <= history_4; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_4 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_4 <= history_5; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_5 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_5 <= history_6; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_6 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_6 <= history_7; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_7 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_7 <= history_8; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_8 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_8 <= history_9; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_9 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_9 <= history_10; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_10 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_10 <= history_11; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_11 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_11 <= history_12; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_12 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_12 <= history_13; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_13 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_13 <= history_14; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_14 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_14 <= history_15; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_15 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_15 <= history_16; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_16 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_16 <= history_17; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_17 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_17 <= history_18; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_18 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_18 <= history_19; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_19 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_19 <= history_20; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_20 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_20 <= history_21; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_21 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_21 <= history_22; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_22 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_22 <= history_23; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_23 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_23 <= history_24; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_24 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_24 <= history_25; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_25 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_25 <= history_26; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_26 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_26 <= history_27; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_27 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_27 <= history_28; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_28 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_28 <= history_29; // @[\\src\\main\\scala\\LFSR.scala 26:16]
    end
    if (reset) begin // @[\\src\\main\\scala\\LFSR.scala 22:24]
      history_29 <= 10'h0; // @[\\src\\main\\scala\\LFSR.scala 22:24]
    end else begin
      history_29 <= {{1'd0}, current_output}; // @[\\src\\main\\scala\\LFSR.scala 28:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_ = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  history_0 = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  history_1 = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  history_2 = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  history_3 = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  history_4 = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  history_5 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  history_6 = _RAND_7[9:0];
  _RAND_8 = {1{`RANDOM}};
  history_7 = _RAND_8[9:0];
  _RAND_9 = {1{`RANDOM}};
  history_8 = _RAND_9[9:0];
  _RAND_10 = {1{`RANDOM}};
  history_9 = _RAND_10[9:0];
  _RAND_11 = {1{`RANDOM}};
  history_10 = _RAND_11[9:0];
  _RAND_12 = {1{`RANDOM}};
  history_11 = _RAND_12[9:0];
  _RAND_13 = {1{`RANDOM}};
  history_12 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  history_13 = _RAND_14[9:0];
  _RAND_15 = {1{`RANDOM}};
  history_14 = _RAND_15[9:0];
  _RAND_16 = {1{`RANDOM}};
  history_15 = _RAND_16[9:0];
  _RAND_17 = {1{`RANDOM}};
  history_16 = _RAND_17[9:0];
  _RAND_18 = {1{`RANDOM}};
  history_17 = _RAND_18[9:0];
  _RAND_19 = {1{`RANDOM}};
  history_18 = _RAND_19[9:0];
  _RAND_20 = {1{`RANDOM}};
  history_19 = _RAND_20[9:0];
  _RAND_21 = {1{`RANDOM}};
  history_20 = _RAND_21[9:0];
  _RAND_22 = {1{`RANDOM}};
  history_21 = _RAND_22[9:0];
  _RAND_23 = {1{`RANDOM}};
  history_22 = _RAND_23[9:0];
  _RAND_24 = {1{`RANDOM}};
  history_23 = _RAND_24[9:0];
  _RAND_25 = {1{`RANDOM}};
  history_24 = _RAND_25[9:0];
  _RAND_26 = {1{`RANDOM}};
  history_25 = _RAND_26[9:0];
  _RAND_27 = {1{`RANDOM}};
  history_26 = _RAND_27[9:0];
  _RAND_28 = {1{`RANDOM}};
  history_27 = _RAND_28[9:0];
  _RAND_29 = {1{`RANDOM}};
  history_28 = _RAND_29[9:0];
  _RAND_30 = {1{`RANDOM}};
  history_29 = _RAND_30[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GameLogic(
  input         clock,
  input         reset,
  input         io_btnC, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnU, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnL, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnR, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_btnD, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_3, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_7, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_8, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_9, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_10, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_11, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_12, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_13, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_14, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_46, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_47, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_48, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_49, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_50, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_51, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_52, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_53, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_54, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_55, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_56, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_57, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_61, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_62, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [10:0] io_spriteXPosition_63, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_3, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_7, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_8, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_9, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_10, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_11, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_12, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_13, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_14, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_46, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_47, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_48, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_49, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_50, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_51, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_52, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_53, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_54, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_55, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_56, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_57, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_61, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_62, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_spriteYPosition_63, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_3, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_4, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_5, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_6, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_7, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_8, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_9, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_10, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_11, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_12, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_13, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_14, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_15, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_46, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_47, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_48, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_49, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_50, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_51, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_52, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_53, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_54, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_55, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_56, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_57, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_61, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_62, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteVisible_63, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpHorizontal_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_16, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_17, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_18, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_19, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_20, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_21, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_22, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_23, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_24, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_25, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_26, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_27, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_28, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_29, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_30, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_31, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_32, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_33, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_34, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_35, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_36, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_37, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_38, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_39, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_40, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_41, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_42, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_43, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_44, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_45, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_58, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_59, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_spriteScaleUpVertical_60, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [9:0]  io_viewBoxX, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output [8:0]  io_viewBoxY, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  input         io_newFrame, // @[\\src\\main\\scala\\GameLogic.scala 12:14]
  output        io_frameUpdateDone // @[\\src\\main\\scala\\GameLogic.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
`endif // RANDOMIZE_REG_INIT
  wire  difficulty_clock; // @[\\src\\main\\scala\\GameLogic.scala 209:26]
  wire  difficulty_reset; // @[\\src\\main\\scala\\GameLogic.scala 209:26]
  wire [1:0] difficulty_io_level; // @[\\src\\main\\scala\\GameLogic.scala 209:26]
  wire [26:0] difficulty_io_speed; // @[\\src\\main\\scala\\GameLogic.scala 209:26]
  wire  difficulty_io_resetSpeed; // @[\\src\\main\\scala\\GameLogic.scala 209:26]
  wire  lfsr_clock; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire  lfsr_reset; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_0; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_1; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_2; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_3; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_4; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_5; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_6; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_7; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_8; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_9; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_10; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_11; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_12; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_13; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_14; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_15; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_16; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_17; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_18; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_19; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_20; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_21; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_22; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_23; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_24; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_25; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_26; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_27; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_28; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  wire [9:0] lfsr_io_out_29; // @[\\src\\main\\scala\\GameLogic.scala 250:20]
  reg [2:0] stateReg; // @[\\src\\main\\scala\\GameLogic.scala 113:25]
  reg [10:0] spriteXRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [10:0] spriteXRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
  reg [9:0] spriteYRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg [9:0] spriteYRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
  reg  spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteVisibleRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
  reg  spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
  reg  initializePositions; // @[\\src\\main\\scala\\GameLogic.scala 130:36]
  wire [10:0] _GEN_0 = initializePositions ? $signed(11'sh140) : $signed(spriteXRegs_3); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_1 = initializePositions ? $signed(10'shf0) : $signed(spriteYRegs_3); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_14 = initializePositions ? $signed(11'sh140) : $signed(spriteXRegs_13); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_15 = initializePositions ? $signed(10'shf0) : $signed(spriteYRegs_13); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_16 = initializePositions ? $signed(11'sh260) : $signed(spriteXRegs_14); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_17 = initializePositions ? $signed(10'shf0) : $signed(spriteYRegs_14); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_18 = initializePositions ? $signed(11'sh168) : $signed(spriteXRegs_16); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_19 = initializePositions ? $signed(10'sh14) : $signed(spriteYRegs_16); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_20 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_17); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_21 = initializePositions ? $signed(10'sh32) : $signed(spriteYRegs_17); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_22 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_18); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_23 = initializePositions ? $signed(10'sh50) : $signed(spriteYRegs_18); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_24 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_19); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_25 = initializePositions ? $signed(10'sh6e) : $signed(spriteYRegs_19); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_26 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_20); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_27 = initializePositions ? $signed(10'sh8c) : $signed(spriteYRegs_20); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_28 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_21); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_29 = initializePositions ? $signed(10'shaa) : $signed(spriteYRegs_21); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_30 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_22); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_31 = initializePositions ? $signed(10'shc8) : $signed(spriteYRegs_22); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_32 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_23); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_33 = initializePositions ? $signed(10'she6) : $signed(spriteYRegs_23); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_34 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_24); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_35 = initializePositions ? $signed(10'sh104) : $signed(spriteYRegs_24); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_36 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_25); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_37 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_25); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_38 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_26); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_39 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_26); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_40 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_27); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_41 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_27); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_42 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_28); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_43 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_28); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_44 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_29); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_45 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_29); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_46 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_30); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_47 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_30); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_48 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_31); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_49 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_31); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_50 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_32); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_51 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_32); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_52 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_33); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_53 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_33); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_54 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_34); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_55 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_34); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_56 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_35); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_57 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_35); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_58 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_36); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_59 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_36); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_60 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_37); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_61 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_37); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_62 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_38); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_63 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_38); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_64 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_39); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_65 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_39); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_66 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_40); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_67 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_40); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_68 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_41); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_69 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_41); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_70 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_42); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_71 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_42); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_72 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_43); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_73 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_43); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_74 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_44); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_75 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_44); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_76 = initializePositions ? $signed(11'sh14) : $signed(spriteXRegs_45); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_77 = initializePositions ? $signed(10'sh122) : $signed(spriteYRegs_45); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_102 = initializePositions ? $signed(11'sh140) : $signed(spriteXRegs_58); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_103 = initializePositions ? $signed(10'sh14) : $signed(spriteYRegs_58); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_104 = initializePositions ? $signed(11'sh1f4) : $signed(spriteXRegs_59); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_105 = initializePositions ? $signed(10'sh46) : $signed(spriteYRegs_59); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire [10:0] _GEN_106 = initializePositions ? $signed(11'sh96) : $signed(spriteXRegs_60); // @[\\src\\main\\scala\\GameLogic.scala 131:29 161:23 121:28]
  wire [9:0] _GEN_107 = initializePositions ? $signed(10'sh64) : $signed(spriteYRegs_60); // @[\\src\\main\\scala\\GameLogic.scala 131:29 162:23 122:28]
  wire  _GEN_114 = initializePositions ? 1'h0 : initializePositions; // @[\\src\\main\\scala\\GameLogic.scala 131:29 164:25 130:36]
  reg  sprite58ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 168:42]
  reg  sprite58ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 169:40]
  reg  sprite59ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 170:42]
  reg  sprite59ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 171:40]
  reg  sprite60ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 172:42]
  reg  sprite60ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 173:40]
  reg [9:0] viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 201:28]
  reg [8:0] viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 202:28]
  reg [1:0] lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 211:23]
  reg [2:0] livesReg; // @[\\src\\main\\scala\\GameLogic.scala 222:25]
  reg [9:0] extraLifeCnt; // @[\\src\\main\\scala\\GameLogic.scala 225:29]
  wire  _difficulty_io_resetSpeed_T_1 = livesReg == 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 228:62]
  reg [7:0] spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 231:34]
  reg [5:0] nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 232:34]
  reg [9:0] starCnt; // @[\\src\\main\\scala\\GameLogic.scala 235:24]
  reg  collisionDetected; // @[\\src\\main\\scala\\GameLogic.scala 238:34]
  reg [7:0] blinkCounter; // @[\\src\\main\\scala\\GameLogic.scala 239:29]
  reg [1:0] blinkTimes; // @[\\src\\main\\scala\\GameLogic.scala 240:27]
  reg  isBlinking; // @[\\src\\main\\scala\\GameLogic.scala 241:27]
  reg  gameOverReturnPressed; // @[\\src\\main\\scala\\GameLogic.scala 247:38]
  wire  _T = lvlReg != 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 253:15]
  wire  _T_2 = livesReg == 3'h2; // @[\\src\\main\\scala\\GameLogic.scala 258:25]
  wire  _T_3 = livesReg == 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 262:25]
  wire  _GEN_117 = livesReg == 3'h2 | _T_3; // @[\\src\\main\\scala\\GameLogic.scala 258:34 259:29]
  wire  _GEN_120 = _difficulty_io_resetSpeed_T_1 | _GEN_117; // @[\\src\\main\\scala\\GameLogic.scala 254:28 255:29]
  wire  _GEN_121 = _difficulty_io_resetSpeed_T_1 | _T_2; // @[\\src\\main\\scala\\GameLogic.scala 254:28 256:29]
  wire  _GEN_123 = lvlReg != 2'h0 & _GEN_120; // @[\\src\\main\\scala\\GameLogic.scala 253:24 272:27]
  wire  _GEN_124 = lvlReg != 2'h0 & _GEN_121; // @[\\src\\main\\scala\\GameLogic.scala 253:24 273:27]
  wire  _GEN_125 = lvlReg != 2'h0 & _difficulty_io_resetSpeed_T_1; // @[\\src\\main\\scala\\GameLogic.scala 253:24 274:27]
  wire  _T_5 = livesReg == 3'h0; // @[\\src\\main\\scala\\GameLogic.scala 343:29]
  wire [2:0] _GEN_126 = livesReg == 3'h0 ? 3'h6 : 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 343:38 344:20 346:20]
  wire  _GEN_138 = gameOverReturnPressed | _GEN_114; // @[\\src\\main\\scala\\GameLogic.scala 293:25 339:37]
  wire  _GEN_139 = gameOverReturnPressed | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 296:26 125:34 339:37]
  wire  _GEN_196 = io_newFrame ? _GEN_138 : _GEN_114; // @[\\src\\main\\scala\\GameLogic.scala 338:25]
  wire [9:0] _spriteYRegs_16_T_2 = 10'h64 + lfsr_io_out_0; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_129 = {{16{spriteXRegs_16[10]}},spriteXRegs_16}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_16_T_2 = $signed(_GEN_129) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_243 = spriteVisibleRegs_16 ? $signed(_spriteXRegs_16_T_2) : $signed({{16{_GEN_18[10]}},_GEN_18}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_244 = $signed(spriteXRegs_16) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_243); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_245 = $signed(spriteXRegs_16) >= 11'sh280 ? $signed(_spriteYRegs_16_T_2) : $signed(_GEN_19); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_246 = $signed(spriteXRegs_16) >= 11'sh280 ? lfsr_io_out_10[0] : spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_247 = ~spriteScaleTypeRegs_0 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [9:0] _spriteYRegs_17_T_2 = 10'h64 + lfsr_io_out_1; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_187 = {{16{spriteXRegs_17[10]}},spriteXRegs_17}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_17_T_2 = $signed(_GEN_187) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_248 = spriteVisibleRegs_17 ? $signed(_spriteXRegs_17_T_2) : $signed({{16{_GEN_20[10]}},_GEN_20}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_249 = $signed(spriteXRegs_17) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_248); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_250 = $signed(spriteXRegs_17) >= 11'sh280 ? $signed(_spriteYRegs_17_T_2) : $signed(_GEN_21); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_251 = $signed(spriteXRegs_17) >= 11'sh280 ? lfsr_io_out_11[0] : spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_252 = ~spriteScaleTypeRegs_1 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [9:0] _spriteYRegs_18_T_2 = 10'h64 + lfsr_io_out_2; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_533 = {{16{spriteXRegs_18[10]}},spriteXRegs_18}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_18_T_2 = $signed(_GEN_533) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_253 = spriteVisibleRegs_18 ? $signed(_spriteXRegs_18_T_2) : $signed({{16{_GEN_22[10]}},_GEN_22}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_254 = $signed(spriteXRegs_18) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_253); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_255 = $signed(spriteXRegs_18) >= 11'sh280 ? $signed(_spriteYRegs_18_T_2) : $signed(_GEN_23); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_256 = $signed(spriteXRegs_18) >= 11'sh280 ? lfsr_io_out_12[0] : spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_257 = ~spriteScaleTypeRegs_2 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [9:0] _spriteYRegs_19_T_2 = 10'h64 + lfsr_io_out_3; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_534 = {{16{spriteXRegs_19[10]}},spriteXRegs_19}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_19_T_2 = $signed(_GEN_534) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_258 = spriteVisibleRegs_19 ? $signed(_spriteXRegs_19_T_2) : $signed({{16{_GEN_24[10]}},_GEN_24}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_259 = $signed(spriteXRegs_19) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_258); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_260 = $signed(spriteXRegs_19) >= 11'sh280 ? $signed(_spriteYRegs_19_T_2) : $signed(_GEN_25); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_261 = $signed(spriteXRegs_19) >= 11'sh280 ? lfsr_io_out_13[0] : spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_262 = ~spriteScaleTypeRegs_3 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [9:0] _spriteYRegs_20_T_2 = 10'h64 + lfsr_io_out_4; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_535 = {{16{spriteXRegs_20[10]}},spriteXRegs_20}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_20_T_2 = $signed(_GEN_535) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_263 = spriteVisibleRegs_20 ? $signed(_spriteXRegs_20_T_2) : $signed({{16{_GEN_26[10]}},_GEN_26}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_264 = $signed(spriteXRegs_20) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_263); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_265 = $signed(spriteXRegs_20) >= 11'sh280 ? $signed(_spriteYRegs_20_T_2) : $signed(_GEN_27); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_266 = $signed(spriteXRegs_20) >= 11'sh280 ? lfsr_io_out_14[0] : spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_267 = ~spriteScaleTypeRegs_4 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [9:0] _spriteYRegs_21_T_2 = 10'h64 + lfsr_io_out_5; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_591 = {{16{spriteXRegs_21[10]}},spriteXRegs_21}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_21_T_2 = $signed(_GEN_591) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_268 = spriteVisibleRegs_21 ? $signed(_spriteXRegs_21_T_2) : $signed({{16{_GEN_28[10]}},_GEN_28}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_269 = $signed(spriteXRegs_21) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_268); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_270 = $signed(spriteXRegs_21) >= 11'sh280 ? $signed(_spriteYRegs_21_T_2) : $signed(_GEN_29); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_271 = $signed(spriteXRegs_21) >= 11'sh280 ? lfsr_io_out_15[0] : spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_272 = ~spriteScaleTypeRegs_5 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [9:0] _spriteYRegs_22_T_2 = 10'h64 + lfsr_io_out_6; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_592 = {{16{spriteXRegs_22[10]}},spriteXRegs_22}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_22_T_2 = $signed(_GEN_592) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_273 = spriteVisibleRegs_22 ? $signed(_spriteXRegs_22_T_2) : $signed({{16{_GEN_30[10]}},_GEN_30}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_274 = $signed(spriteXRegs_22) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_273); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_275 = $signed(spriteXRegs_22) >= 11'sh280 ? $signed(_spriteYRegs_22_T_2) : $signed(_GEN_31); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_276 = $signed(spriteXRegs_22) >= 11'sh280 ? lfsr_io_out_16[0] : spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_277 = ~spriteScaleTypeRegs_6 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [9:0] _spriteYRegs_23_T_2 = 10'h64 + lfsr_io_out_7; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_593 = {{16{spriteXRegs_23[10]}},spriteXRegs_23}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_23_T_2 = $signed(_GEN_593) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_278 = spriteVisibleRegs_23 ? $signed(_spriteXRegs_23_T_2) : $signed({{16{_GEN_32[10]}},_GEN_32}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_279 = $signed(spriteXRegs_23) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_278); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_280 = $signed(spriteXRegs_23) >= 11'sh280 ? $signed(_spriteYRegs_23_T_2) : $signed(_GEN_33); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_281 = $signed(spriteXRegs_23) >= 11'sh280 ? lfsr_io_out_17[0] : spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_282 = ~spriteScaleTypeRegs_7 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [9:0] _spriteYRegs_24_T_2 = 10'h64 + lfsr_io_out_8; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_598 = {{16{spriteXRegs_24[10]}},spriteXRegs_24}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_24_T_2 = $signed(_GEN_598) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_283 = spriteVisibleRegs_24 ? $signed(_spriteXRegs_24_T_2) : $signed({{16{_GEN_34[10]}},_GEN_34}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_284 = $signed(spriteXRegs_24) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_283); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_285 = $signed(spriteXRegs_24) >= 11'sh280 ? $signed(_spriteYRegs_24_T_2) : $signed(_GEN_35); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_286 = $signed(spriteXRegs_24) >= 11'sh280 ? lfsr_io_out_18[0] : spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_287 = ~spriteScaleTypeRegs_8 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [9:0] _spriteYRegs_25_T_2 = 10'h64 + lfsr_io_out_9; // @[\\src\\main\\scala\\GameLogic.scala 367:63]
  wire [26:0] _GEN_599 = {{16{spriteXRegs_25[10]}},spriteXRegs_25}; // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _spriteXRegs_25_T_2 = $signed(_GEN_599) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 372:46]
  wire [26:0] _GEN_288 = spriteVisibleRegs_25 ? $signed(_spriteXRegs_25_T_2) : $signed({{16{_GEN_36[10]}},_GEN_36}); // @[\\src\\main\\scala\\GameLogic.scala 371:44 372:28]
  wire [26:0] _GEN_289 = $signed(spriteXRegs_25) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_288); // @[\\src\\main\\scala\\GameLogic.scala 365:41 366:28]
  wire [9:0] _GEN_290 = $signed(spriteXRegs_25) >= 11'sh280 ? $signed(_spriteYRegs_25_T_2) : $signed(_GEN_37); // @[\\src\\main\\scala\\GameLogic.scala 365:41 367:28]
  wire  _GEN_291 = $signed(spriteXRegs_25) >= 11'sh280 ? lfsr_io_out_19[0] : spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 126:36 365:41 369:40]
  wire  _GEN_292 = ~spriteScaleTypeRegs_9 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 376:52 377:43 380:43]
  wire [26:0] _GEN_600 = {{16{spriteXRegs_26[10]}},spriteXRegs_26}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_26_T_2 = $signed(_GEN_600) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_293 = spriteVisibleRegs_26 ? $signed(_spriteXRegs_26_T_2) : $signed({{16{_GEN_38[10]}},_GEN_38}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_294 = $signed(spriteXRegs_26) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_293); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_295 = $signed(spriteXRegs_26) >= 11'sh280 ? $signed(_spriteYRegs_16_T_2) : $signed(_GEN_39); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_296 = $signed(spriteXRegs_26) >= 11'sh280 ? lfsr_io_out_10[0] : _GEN_246; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [26:0] _GEN_656 = {{16{spriteXRegs_27[10]}},spriteXRegs_27}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_27_T_2 = $signed(_GEN_656) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_298 = spriteVisibleRegs_27 ? $signed(_spriteXRegs_27_T_2) : $signed({{16{_GEN_40[10]}},_GEN_40}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_299 = $signed(spriteXRegs_27) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_298); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_300 = $signed(spriteXRegs_27) >= 11'sh280 ? $signed(_spriteYRegs_17_T_2) : $signed(_GEN_41); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_301 = $signed(spriteXRegs_27) >= 11'sh280 ? lfsr_io_out_11[0] : _GEN_251; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [26:0] _GEN_657 = {{16{spriteXRegs_28[10]}},spriteXRegs_28}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_28_T_2 = $signed(_GEN_657) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_303 = spriteVisibleRegs_28 ? $signed(_spriteXRegs_28_T_2) : $signed({{16{_GEN_42[10]}},_GEN_42}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_304 = $signed(spriteXRegs_28) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_303); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_305 = $signed(spriteXRegs_28) >= 11'sh280 ? $signed(_spriteYRegs_18_T_2) : $signed(_GEN_43); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_306 = $signed(spriteXRegs_28) >= 11'sh280 ? lfsr_io_out_12[0] : _GEN_256; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [26:0] _GEN_658 = {{16{spriteXRegs_29[10]}},spriteXRegs_29}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_29_T_2 = $signed(_GEN_658) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_308 = spriteVisibleRegs_29 ? $signed(_spriteXRegs_29_T_2) : $signed({{16{_GEN_44[10]}},_GEN_44}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_309 = $signed(spriteXRegs_29) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_308); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_310 = $signed(spriteXRegs_29) >= 11'sh280 ? $signed(_spriteYRegs_19_T_2) : $signed(_GEN_45); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_311 = $signed(spriteXRegs_29) >= 11'sh280 ? lfsr_io_out_13[0] : _GEN_261; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [26:0] _GEN_664 = {{16{spriteXRegs_30[10]}},spriteXRegs_30}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_30_T_2 = $signed(_GEN_664) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_313 = spriteVisibleRegs_30 ? $signed(_spriteXRegs_30_T_2) : $signed({{16{_GEN_46[10]}},_GEN_46}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_314 = $signed(spriteXRegs_30) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_313); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_315 = $signed(spriteXRegs_30) >= 11'sh280 ? $signed(_spriteYRegs_20_T_2) : $signed(_GEN_47); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_316 = $signed(spriteXRegs_30) >= 11'sh280 ? lfsr_io_out_14[0] : _GEN_266; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [26:0] _GEN_665 = {{16{spriteXRegs_31[10]}},spriteXRegs_31}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_31_T_2 = $signed(_GEN_665) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_318 = spriteVisibleRegs_31 ? $signed(_spriteXRegs_31_T_2) : $signed({{16{_GEN_48[10]}},_GEN_48}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_319 = $signed(spriteXRegs_31) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_318); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_320 = $signed(spriteXRegs_31) >= 11'sh280 ? $signed(_spriteYRegs_21_T_2) : $signed(_GEN_49); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_321 = $signed(spriteXRegs_31) >= 11'sh280 ? lfsr_io_out_15[0] : _GEN_271; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [26:0] _GEN_666 = {{16{spriteXRegs_32[10]}},spriteXRegs_32}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_32_T_2 = $signed(_GEN_666) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_323 = spriteVisibleRegs_32 ? $signed(_spriteXRegs_32_T_2) : $signed({{16{_GEN_50[10]}},_GEN_50}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_324 = $signed(spriteXRegs_32) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_323); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_325 = $signed(spriteXRegs_32) >= 11'sh280 ? $signed(_spriteYRegs_22_T_2) : $signed(_GEN_51); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_326 = $signed(spriteXRegs_32) >= 11'sh280 ? lfsr_io_out_16[0] : _GEN_276; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [26:0] _GEN_722 = {{16{spriteXRegs_33[10]}},spriteXRegs_33}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_33_T_2 = $signed(_GEN_722) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_328 = spriteVisibleRegs_33 ? $signed(_spriteXRegs_33_T_2) : $signed({{16{_GEN_52[10]}},_GEN_52}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_329 = $signed(spriteXRegs_33) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_328); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_330 = $signed(spriteXRegs_33) >= 11'sh280 ? $signed(_spriteYRegs_23_T_2) : $signed(_GEN_53); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_331 = $signed(spriteXRegs_33) >= 11'sh280 ? lfsr_io_out_17[0] : _GEN_281; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [26:0] _GEN_723 = {{16{spriteXRegs_34[10]}},spriteXRegs_34}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_34_T_2 = $signed(_GEN_723) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_333 = spriteVisibleRegs_34 ? $signed(_spriteXRegs_34_T_2) : $signed({{16{_GEN_54[10]}},_GEN_54}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_334 = $signed(spriteXRegs_34) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_333); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_335 = $signed(spriteXRegs_34) >= 11'sh280 ? $signed(_spriteYRegs_24_T_2) : $signed(_GEN_55); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_336 = $signed(spriteXRegs_34) >= 11'sh280 ? lfsr_io_out_18[0] : _GEN_286; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [26:0] _GEN_724 = {{16{spriteXRegs_35[10]}},spriteXRegs_35}; // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _spriteXRegs_35_T_2 = $signed(_GEN_724) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 395:46]
  wire [26:0] _GEN_338 = spriteVisibleRegs_35 ? $signed(_spriteXRegs_35_T_2) : $signed({{16{_GEN_56[10]}},_GEN_56}); // @[\\src\\main\\scala\\GameLogic.scala 394:44 395:28]
  wire [26:0] _GEN_339 = $signed(spriteXRegs_35) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_338); // @[\\src\\main\\scala\\GameLogic.scala 388:41 389:28]
  wire [9:0] _GEN_340 = $signed(spriteXRegs_35) >= 11'sh280 ? $signed(_spriteYRegs_25_T_2) : $signed(_GEN_57); // @[\\src\\main\\scala\\GameLogic.scala 388:41 390:28]
  wire  _GEN_341 = $signed(spriteXRegs_35) >= 11'sh280 ? lfsr_io_out_19[0] : _GEN_291; // @[\\src\\main\\scala\\GameLogic.scala 388:41 392:40]
  wire [9:0] _spriteYRegs_36_T_2 = 10'h64 + lfsr_io_out_20; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_729 = {{16{spriteXRegs_36[10]}},spriteXRegs_36}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_36_T_2 = $signed(_GEN_729) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_343 = spriteVisibleRegs_36 ? $signed(_spriteXRegs_36_T_2) : $signed({{16{_GEN_58[10]}},_GEN_58}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_344 = $signed(spriteXRegs_36) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_343); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_345 = $signed(spriteXRegs_36) >= 11'sh280 ? $signed(_spriteYRegs_36_T_2) : $signed(_GEN_59); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_346 = $signed(spriteXRegs_36) >= 11'sh280 ? lfsr_io_out_10[0] : _GEN_296; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _spriteYRegs_37_T_2 = 10'h64 + lfsr_io_out_21; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_730 = {{16{spriteXRegs_37[10]}},spriteXRegs_37}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_37_T_2 = $signed(_GEN_730) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_348 = spriteVisibleRegs_37 ? $signed(_spriteXRegs_37_T_2) : $signed({{16{_GEN_60[10]}},_GEN_60}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_349 = $signed(spriteXRegs_37) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_348); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_350 = $signed(spriteXRegs_37) >= 11'sh280 ? $signed(_spriteYRegs_37_T_2) : $signed(_GEN_61); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_351 = $signed(spriteXRegs_37) >= 11'sh280 ? lfsr_io_out_11[0] : _GEN_301; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _spriteYRegs_38_T_2 = 10'h64 + lfsr_io_out_22; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_731 = {{16{spriteXRegs_38[10]}},spriteXRegs_38}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_38_T_2 = $signed(_GEN_731) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_353 = spriteVisibleRegs_38 ? $signed(_spriteXRegs_38_T_2) : $signed({{16{_GEN_62[10]}},_GEN_62}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_354 = $signed(spriteXRegs_38) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_353); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_355 = $signed(spriteXRegs_38) >= 11'sh280 ? $signed(_spriteYRegs_38_T_2) : $signed(_GEN_63); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_356 = $signed(spriteXRegs_38) >= 11'sh280 ? lfsr_io_out_12[0] : _GEN_306; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _spriteYRegs_39_T_2 = 10'h64 + lfsr_io_out_23; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_787 = {{16{spriteXRegs_39[10]}},spriteXRegs_39}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_39_T_2 = $signed(_GEN_787) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_358 = spriteVisibleRegs_39 ? $signed(_spriteXRegs_39_T_2) : $signed({{16{_GEN_64[10]}},_GEN_64}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_359 = $signed(spriteXRegs_39) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_358); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_360 = $signed(spriteXRegs_39) >= 11'sh280 ? $signed(_spriteYRegs_39_T_2) : $signed(_GEN_65); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_361 = $signed(spriteXRegs_39) >= 11'sh280 ? lfsr_io_out_13[0] : _GEN_311; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _spriteYRegs_40_T_2 = 10'h64 + lfsr_io_out_24; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_788 = {{16{spriteXRegs_40[10]}},spriteXRegs_40}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_40_T_2 = $signed(_GEN_788) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_363 = spriteVisibleRegs_40 ? $signed(_spriteXRegs_40_T_2) : $signed({{16{_GEN_66[10]}},_GEN_66}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_364 = $signed(spriteXRegs_40) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_363); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_365 = $signed(spriteXRegs_40) >= 11'sh280 ? $signed(_spriteYRegs_40_T_2) : $signed(_GEN_67); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_366 = $signed(spriteXRegs_40) >= 11'sh280 ? lfsr_io_out_14[0] : _GEN_316; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _spriteYRegs_41_T_2 = 10'h64 + lfsr_io_out_25; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_789 = {{16{spriteXRegs_41[10]}},spriteXRegs_41}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_41_T_2 = $signed(_GEN_789) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_368 = spriteVisibleRegs_41 ? $signed(_spriteXRegs_41_T_2) : $signed({{16{_GEN_68[10]}},_GEN_68}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_369 = $signed(spriteXRegs_41) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_368); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_370 = $signed(spriteXRegs_41) >= 11'sh280 ? $signed(_spriteYRegs_41_T_2) : $signed(_GEN_69); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_371 = $signed(spriteXRegs_41) >= 11'sh280 ? lfsr_io_out_15[0] : _GEN_321; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _spriteYRegs_42_T_2 = 10'h64 + lfsr_io_out_26; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_795 = {{16{spriteXRegs_42[10]}},spriteXRegs_42}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_42_T_2 = $signed(_GEN_795) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_373 = spriteVisibleRegs_42 ? $signed(_spriteXRegs_42_T_2) : $signed({{16{_GEN_70[10]}},_GEN_70}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_374 = $signed(spriteXRegs_42) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_373); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_375 = $signed(spriteXRegs_42) >= 11'sh280 ? $signed(_spriteYRegs_42_T_2) : $signed(_GEN_71); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_376 = $signed(spriteXRegs_42) >= 11'sh280 ? lfsr_io_out_16[0] : _GEN_326; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _spriteYRegs_43_T_2 = 10'h64 + lfsr_io_out_27; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_796 = {{16{spriteXRegs_43[10]}},spriteXRegs_43}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_43_T_2 = $signed(_GEN_796) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_378 = spriteVisibleRegs_43 ? $signed(_spriteXRegs_43_T_2) : $signed({{16{_GEN_72[10]}},_GEN_72}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_379 = $signed(spriteXRegs_43) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_378); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_380 = $signed(spriteXRegs_43) >= 11'sh280 ? $signed(_spriteYRegs_43_T_2) : $signed(_GEN_73); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_381 = $signed(spriteXRegs_43) >= 11'sh280 ? lfsr_io_out_17[0] : _GEN_331; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _spriteYRegs_44_T_2 = 10'h64 + lfsr_io_out_28; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_797 = {{16{spriteXRegs_44[10]}},spriteXRegs_44}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_44_T_2 = $signed(_GEN_797) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_383 = spriteVisibleRegs_44 ? $signed(_spriteXRegs_44_T_2) : $signed({{16{_GEN_74[10]}},_GEN_74}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_384 = $signed(spriteXRegs_44) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_383); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_385 = $signed(spriteXRegs_44) >= 11'sh280 ? $signed(_spriteYRegs_44_T_2) : $signed(_GEN_75); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_386 = $signed(spriteXRegs_44) >= 11'sh280 ? lfsr_io_out_18[0] : _GEN_336; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _spriteYRegs_45_T_2 = 10'h64 + lfsr_io_out_29; // @[\\src\\main\\scala\\GameLogic.scala 413:63]
  wire [26:0] _GEN_853 = {{16{spriteXRegs_45[10]}},spriteXRegs_45}; // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _spriteXRegs_45_T_2 = $signed(_GEN_853) + $signed(difficulty_io_speed); // @[\\src\\main\\scala\\GameLogic.scala 419:46]
  wire [26:0] _GEN_388 = spriteVisibleRegs_45 ? $signed(_spriteXRegs_45_T_2) : $signed({{16{_GEN_76[10]}},_GEN_76}); // @[\\src\\main\\scala\\GameLogic.scala 418:44 419:28]
  wire [26:0] _GEN_389 = $signed(spriteXRegs_45) >= 11'sh280 ? $signed(-27'sh20) : $signed(_GEN_388); // @[\\src\\main\\scala\\GameLogic.scala 411:41 412:28]
  wire [9:0] _GEN_390 = $signed(spriteXRegs_45) >= 11'sh280 ? $signed(_spriteYRegs_45_T_2) : $signed(_GEN_77); // @[\\src\\main\\scala\\GameLogic.scala 411:41 413:28]
  wire  _GEN_391 = $signed(spriteXRegs_45) >= 11'sh280 ? lfsr_io_out_19[0] : _GEN_341; // @[\\src\\main\\scala\\GameLogic.scala 411:41 416:40]
  wire [9:0] _extraLifeCnt_T_1 = extraLifeCnt + 10'h1; // @[\\src\\main\\scala\\GameLogic.scala 439:40]
  wire [10:0] _GEN_393 = extraLifeCnt == 10'h258 ? $signed(-11'sh20) : $signed(_GEN_14); // @[\\src\\main\\scala\\GameLogic.scala 433:38 434:27]
  wire  _GEN_394 = extraLifeCnt == 10'h258 | spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 433:38 435:33 125:34]
  wire [9:0] _GEN_395 = extraLifeCnt == 10'h258 ? $signed(lfsr_io_out_0) : $signed(_GEN_15); // @[\\src\\main\\scala\\GameLogic.scala 433:38 436:27]
  wire [9:0] _GEN_396 = extraLifeCnt == 10'h258 ? 10'h0 : _extraLifeCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 433:38 437:24 439:24]
  wire [10:0] _spriteXRegs_13_T_2 = $signed(spriteXRegs_13) + 11'sh2; // @[\\src\\main\\scala\\GameLogic.scala 442:46]
  wire [10:0] _GEN_397 = spriteVisibleRegs_13 ? $signed(_spriteXRegs_13_T_2) : $signed(_GEN_393); // @[\\src\\main\\scala\\GameLogic.scala 441:37 442:27]
  wire  _GEN_398 = $signed(spriteXRegs_13) >= 11'sh280 ? 1'h0 : _GEN_394; // @[\\src\\main\\scala\\GameLogic.scala 444:40 445:33]
  wire [26:0] _GEN_399 = _T ? $signed(_GEN_244) : $signed({{16{_GEN_18[10]}},_GEN_18}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_402 = _T ? _GEN_247 : spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_404 = _T ? $signed(_GEN_249) : $signed({{16{_GEN_20[10]}},_GEN_20}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_407 = _T ? _GEN_252 : spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_409 = _T ? $signed(_GEN_254) : $signed({{16{_GEN_22[10]}},_GEN_22}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_412 = _T ? _GEN_257 : spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_414 = _T ? $signed(_GEN_259) : $signed({{16{_GEN_24[10]}},_GEN_24}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_417 = _T ? _GEN_262 : spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_419 = _T ? $signed(_GEN_264) : $signed({{16{_GEN_26[10]}},_GEN_26}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_422 = _T ? _GEN_267 : spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_424 = _T ? $signed(_GEN_269) : $signed({{16{_GEN_28[10]}},_GEN_28}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_427 = _T ? _GEN_272 : spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_429 = _T ? $signed(_GEN_274) : $signed({{16{_GEN_30[10]}},_GEN_30}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_432 = _T ? _GEN_277 : spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_434 = _T ? $signed(_GEN_279) : $signed({{16{_GEN_32[10]}},_GEN_32}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_437 = _T ? _GEN_282 : spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_439 = _T ? $signed(_GEN_284) : $signed({{16{_GEN_34[10]}},_GEN_34}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_442 = _T ? _GEN_287 : spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_444 = _T ? $signed(_GEN_289) : $signed({{16{_GEN_36[10]}},_GEN_36}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_447 = _T ? _GEN_292 : spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 359:29 187:35]
  wire [26:0] _GEN_449 = _T ? $signed(_GEN_294) : $signed({{16{_GEN_38[10]}},_GEN_38}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_453 = _T ? $signed(_GEN_299) : $signed({{16{_GEN_40[10]}},_GEN_40}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_457 = _T ? $signed(_GEN_304) : $signed({{16{_GEN_42[10]}},_GEN_42}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_461 = _T ? $signed(_GEN_309) : $signed({{16{_GEN_44[10]}},_GEN_44}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_465 = _T ? $signed(_GEN_314) : $signed({{16{_GEN_46[10]}},_GEN_46}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_469 = _T ? $signed(_GEN_319) : $signed({{16{_GEN_48[10]}},_GEN_48}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_473 = _T ? $signed(_GEN_324) : $signed({{16{_GEN_50[10]}},_GEN_50}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_477 = _T ? $signed(_GEN_329) : $signed({{16{_GEN_52[10]}},_GEN_52}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_481 = _T ? $signed(_GEN_334) : $signed({{16{_GEN_54[10]}},_GEN_54}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_485 = _T ? $signed(_GEN_339) : $signed({{16{_GEN_56[10]}},_GEN_56}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_489 = _T ? $signed(_GEN_344) : $signed({{16{_GEN_58[10]}},_GEN_58}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_493 = _T ? $signed(_GEN_349) : $signed({{16{_GEN_60[10]}},_GEN_60}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_497 = _T ? $signed(_GEN_354) : $signed({{16{_GEN_62[10]}},_GEN_62}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_501 = _T ? $signed(_GEN_359) : $signed({{16{_GEN_64[10]}},_GEN_64}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_505 = _T ? $signed(_GEN_364) : $signed({{16{_GEN_66[10]}},_GEN_66}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_509 = _T ? $signed(_GEN_369) : $signed({{16{_GEN_68[10]}},_GEN_68}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_513 = _T ? $signed(_GEN_374) : $signed({{16{_GEN_70[10]}},_GEN_70}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_517 = _T ? $signed(_GEN_379) : $signed({{16{_GEN_72[10]}},_GEN_72}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_521 = _T ? $signed(_GEN_384) : $signed({{16{_GEN_74[10]}},_GEN_74}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire [26:0] _GEN_525 = _T ? $signed(_GEN_389) : $signed({{16{_GEN_76[10]}},_GEN_76}); // @[\\src\\main\\scala\\GameLogic.scala 359:29]
  wire  _GEN_530 = _T ? _GEN_398 : spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 359:29 125:34]
  wire  _T_69 = lvlReg == 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 450:19]
  wire  _T_72 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha; // @[\\src\\main\\scala\\GameLogic.scala 452:40]
  wire [5:0] _T_74 = 6'h10 + nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 453:34]
  wire  _GEN_536 = 6'h3 == _T_74 | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_537 = 6'h4 == _T_74 | spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_538 = 6'h5 == _T_74 | spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_539 = 6'h6 == _T_74 | spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_540 = 6'h7 == _T_74 | spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_541 = 6'h8 == _T_74 | spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_542 = 6'h9 == _T_74 | spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_543 = 6'ha == _T_74 | spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_544 = 6'hb == _T_74 | spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_545 = 6'hc == _T_74 | spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_546 = 6'hd == _T_74 | _GEN_530; // @[\\src\\main\\scala\\GameLogic.scala 453:{55,55}]
  wire  _GEN_547 = 6'he == _T_74 | spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_548 = 6'hf == _T_74 | spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_549 = 6'h10 == _T_74 | spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_550 = 6'h11 == _T_74 | spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_551 = 6'h12 == _T_74 | spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_552 = 6'h13 == _T_74 | spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_553 = 6'h14 == _T_74 | spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_554 = 6'h15 == _T_74 | spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_555 = 6'h16 == _T_74 | spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_556 = 6'h17 == _T_74 | spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_557 = 6'h18 == _T_74 | spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_558 = 6'h19 == _T_74 | spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_559 = 6'h1a == _T_74 | spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_560 = 6'h1b == _T_74 | spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_561 = 6'h1c == _T_74 | spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_562 = 6'h1d == _T_74 | spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_563 = 6'h1e == _T_74 | spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_564 = 6'h1f == _T_74 | spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_565 = 6'h20 == _T_74 | spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_566 = 6'h21 == _T_74 | spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_567 = 6'h22 == _T_74 | spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_568 = 6'h23 == _T_74 | spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_569 = 6'h24 == _T_74 | spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_570 = 6'h25 == _T_74 | spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_571 = 6'h26 == _T_74 | spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_572 = 6'h27 == _T_74 | spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_573 = 6'h28 == _T_74 | spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_574 = 6'h29 == _T_74 | spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_575 = 6'h2a == _T_74 | spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_576 = 6'h2b == _T_74 | spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_577 = 6'h2c == _T_74 | spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_578 = 6'h2d == _T_74 | spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_579 = 6'h2e == _T_74 | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_580 = 6'h2f == _T_74 | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_581 = 6'h30 == _T_74 | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_582 = 6'h31 == _T_74 | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_583 = 6'h32 == _T_74 | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_584 = 6'h33 == _T_74 | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_585 = 6'h34 == _T_74 | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_586 = 6'h35 == _T_74 | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_587 = 6'h36 == _T_74 | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_588 = 6'h37 == _T_74 | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_589 = 6'h38 == _T_74 | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_590 = 6'h39 == _T_74 | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 453:{55,55}]
  wire  _GEN_594 = 6'h3d == _T_74 | _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 453:{55,55}]
  wire  _GEN_595 = 6'h3e == _T_74 | _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 453:{55,55}]
  wire  _GEN_596 = 6'h3f == _T_74 | _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 453:{55,55}]
  wire [5:0] _nextSpriteToSpawn_T_1 = nextSpriteToSpawn + 6'h1; // @[\\src\\main\\scala\\GameLogic.scala 454:50]
  wire [7:0] _spawnDelayCounter_T_1 = spawnDelayCounter - 8'h1; // @[\\src\\main\\scala\\GameLogic.scala 457:50]
  wire [7:0] _GEN_597 = spawnDelayCounter > 8'h0 ? _spawnDelayCounter_T_1 : spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 456:45 457:29 231:34]
  wire  _GEN_601 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_536 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_602 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_537 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_603 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_538 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_604 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_539 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_605 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_540 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_606 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_541 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_607 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_542 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_608 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_543 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_609 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_544 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_610 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_545 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_611 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_546 : _GEN_530; // @[\\src\\main\\scala\\GameLogic.scala 452:69]
  wire  _GEN_612 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_547 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_613 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_548 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_614 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_549 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_615 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_550 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_616 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_551 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_617 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_552 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_618 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_553 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_619 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_554 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_620 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_555 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_621 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_556 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_622 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_557 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_623 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_558 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_624 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_559 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_625 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_560 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_626 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_561 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_627 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_562 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_628 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_563 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_629 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_564 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_630 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_565 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_631 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_566 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_632 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_567 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_633 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_568 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_634 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_569 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_635 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_570 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_636 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_571 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_637 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_572 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_638 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_573 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_639 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_574 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_640 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_575 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_641 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_576 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_642 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_577 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_643 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_578 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_644 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_579 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_645 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_580 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_646 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_581 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_647 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_582 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_648 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_583 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_649 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_584 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_650 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_585 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_651 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_586 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_652 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_587 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_653 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_588 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_654 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_589 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_655 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_590 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 452:69]
  wire  _GEN_659 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_594 : _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 452:69]
  wire  _GEN_660 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_595 : _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 452:69]
  wire  _GEN_661 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _GEN_596 : _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 452:69]
  wire [5:0] _GEN_662 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? _nextSpriteToSpawn_T_1 :
    nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 452:69 454:29 232:34]
  wire [7:0] _GEN_663 = spawnDelayCounter == 8'h0 & nextSpriteToSpawn < 6'ha ? 8'h1e : _GEN_597; // @[\\src\\main\\scala\\GameLogic.scala 452:69 455:29]
  wire  _T_76 = lvlReg == 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 459:25]
  wire [5:0] _T_81 = 6'h1a + nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 462:34]
  wire  _GEN_667 = 6'h3 == _T_81 | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_668 = 6'h4 == _T_81 | spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_669 = 6'h5 == _T_81 | spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_670 = 6'h6 == _T_81 | spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_671 = 6'h7 == _T_81 | spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_672 = 6'h8 == _T_81 | spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_673 = 6'h9 == _T_81 | spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_674 = 6'ha == _T_81 | spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_675 = 6'hb == _T_81 | spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_676 = 6'hc == _T_81 | spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_677 = 6'hd == _T_81 | _GEN_530; // @[\\src\\main\\scala\\GameLogic.scala 462:{55,55}]
  wire  _GEN_678 = 6'he == _T_81 | spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_679 = 6'hf == _T_81 | spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_680 = 6'h10 == _T_81 | spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_681 = 6'h11 == _T_81 | spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_682 = 6'h12 == _T_81 | spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_683 = 6'h13 == _T_81 | spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_684 = 6'h14 == _T_81 | spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_685 = 6'h15 == _T_81 | spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_686 = 6'h16 == _T_81 | spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_687 = 6'h17 == _T_81 | spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_688 = 6'h18 == _T_81 | spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_689 = 6'h19 == _T_81 | spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_690 = 6'h1a == _T_81 | spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_691 = 6'h1b == _T_81 | spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_692 = 6'h1c == _T_81 | spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_693 = 6'h1d == _T_81 | spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_694 = 6'h1e == _T_81 | spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_695 = 6'h1f == _T_81 | spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_696 = 6'h20 == _T_81 | spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_697 = 6'h21 == _T_81 | spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_698 = 6'h22 == _T_81 | spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_699 = 6'h23 == _T_81 | spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_700 = 6'h24 == _T_81 | spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_701 = 6'h25 == _T_81 | spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_702 = 6'h26 == _T_81 | spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_703 = 6'h27 == _T_81 | spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_704 = 6'h28 == _T_81 | spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_705 = 6'h29 == _T_81 | spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_706 = 6'h2a == _T_81 | spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_707 = 6'h2b == _T_81 | spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_708 = 6'h2c == _T_81 | spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_709 = 6'h2d == _T_81 | spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_710 = 6'h2e == _T_81 | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_711 = 6'h2f == _T_81 | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_712 = 6'h30 == _T_81 | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_713 = 6'h31 == _T_81 | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_714 = 6'h32 == _T_81 | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_715 = 6'h33 == _T_81 | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_716 = 6'h34 == _T_81 | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_717 = 6'h35 == _T_81 | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_718 = 6'h36 == _T_81 | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_719 = 6'h37 == _T_81 | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_720 = 6'h38 == _T_81 | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_721 = 6'h39 == _T_81 | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 462:{55,55}]
  wire  _GEN_725 = 6'h3d == _T_81 | _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 462:{55,55}]
  wire  _GEN_726 = 6'h3e == _T_81 | _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 462:{55,55}]
  wire  _GEN_727 = 6'h3f == _T_81 | _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 462:{55,55}]
  wire  _GEN_732 = _T_72 ? _GEN_667 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_733 = _T_72 ? _GEN_668 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_734 = _T_72 ? _GEN_669 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_735 = _T_72 ? _GEN_670 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_736 = _T_72 ? _GEN_671 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_737 = _T_72 ? _GEN_672 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_738 = _T_72 ? _GEN_673 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_739 = _T_72 ? _GEN_674 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_740 = _T_72 ? _GEN_675 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_741 = _T_72 ? _GEN_676 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_742 = _T_72 ? _GEN_677 : _GEN_530; // @[\\src\\main\\scala\\GameLogic.scala 461:69]
  wire  _GEN_743 = _T_72 ? _GEN_678 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_744 = _T_72 ? _GEN_679 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_745 = _T_72 ? _GEN_680 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_746 = _T_72 ? _GEN_681 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_747 = _T_72 ? _GEN_682 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_748 = _T_72 ? _GEN_683 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_749 = _T_72 ? _GEN_684 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_750 = _T_72 ? _GEN_685 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_751 = _T_72 ? _GEN_686 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_752 = _T_72 ? _GEN_687 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_753 = _T_72 ? _GEN_688 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_754 = _T_72 ? _GEN_689 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_755 = _T_72 ? _GEN_690 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_756 = _T_72 ? _GEN_691 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_757 = _T_72 ? _GEN_692 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_758 = _T_72 ? _GEN_693 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_759 = _T_72 ? _GEN_694 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_760 = _T_72 ? _GEN_695 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_761 = _T_72 ? _GEN_696 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_762 = _T_72 ? _GEN_697 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_763 = _T_72 ? _GEN_698 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_764 = _T_72 ? _GEN_699 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_765 = _T_72 ? _GEN_700 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_766 = _T_72 ? _GEN_701 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_767 = _T_72 ? _GEN_702 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_768 = _T_72 ? _GEN_703 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_769 = _T_72 ? _GEN_704 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_770 = _T_72 ? _GEN_705 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_771 = _T_72 ? _GEN_706 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_772 = _T_72 ? _GEN_707 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_773 = _T_72 ? _GEN_708 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_774 = _T_72 ? _GEN_709 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_775 = _T_72 ? _GEN_710 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_776 = _T_72 ? _GEN_711 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_777 = _T_72 ? _GEN_712 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_778 = _T_72 ? _GEN_713 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_779 = _T_72 ? _GEN_714 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_780 = _T_72 ? _GEN_715 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_781 = _T_72 ? _GEN_716 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_782 = _T_72 ? _GEN_717 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_783 = _T_72 ? _GEN_718 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_784 = _T_72 ? _GEN_719 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_785 = _T_72 ? _GEN_720 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_786 = _T_72 ? _GEN_721 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 461:69]
  wire  _GEN_790 = _T_72 ? _GEN_725 : _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 461:69]
  wire  _GEN_791 = _T_72 ? _GEN_726 : _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 461:69]
  wire  _GEN_792 = _T_72 ? _GEN_727 : _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 461:69]
  wire [7:0] _GEN_794 = _T_72 ? 8'h19 : _GEN_597; // @[\\src\\main\\scala\\GameLogic.scala 461:69 464:29]
  wire  _T_83 = lvlReg == 2'h3; // @[\\src\\main\\scala\\GameLogic.scala 468:25]
  wire [5:0] _T_88 = 6'h24 + nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 471:34]
  wire  _GEN_798 = 6'h3 == _T_88 | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_799 = 6'h4 == _T_88 | spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_800 = 6'h5 == _T_88 | spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_801 = 6'h6 == _T_88 | spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_802 = 6'h7 == _T_88 | spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_803 = 6'h8 == _T_88 | spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_804 = 6'h9 == _T_88 | spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_805 = 6'ha == _T_88 | spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_806 = 6'hb == _T_88 | spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_807 = 6'hc == _T_88 | spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_808 = 6'hd == _T_88 | _GEN_530; // @[\\src\\main\\scala\\GameLogic.scala 471:{55,55}]
  wire  _GEN_809 = 6'he == _T_88 | spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_810 = 6'hf == _T_88 | spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_811 = 6'h10 == _T_88 | spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_812 = 6'h11 == _T_88 | spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_813 = 6'h12 == _T_88 | spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_814 = 6'h13 == _T_88 | spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_815 = 6'h14 == _T_88 | spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_816 = 6'h15 == _T_88 | spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_817 = 6'h16 == _T_88 | spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_818 = 6'h17 == _T_88 | spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_819 = 6'h18 == _T_88 | spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_820 = 6'h19 == _T_88 | spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_821 = 6'h1a == _T_88 | spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_822 = 6'h1b == _T_88 | spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_823 = 6'h1c == _T_88 | spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_824 = 6'h1d == _T_88 | spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_825 = 6'h1e == _T_88 | spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_826 = 6'h1f == _T_88 | spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_827 = 6'h20 == _T_88 | spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_828 = 6'h21 == _T_88 | spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_829 = 6'h22 == _T_88 | spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_830 = 6'h23 == _T_88 | spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_831 = 6'h24 == _T_88 | spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_832 = 6'h25 == _T_88 | spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_833 = 6'h26 == _T_88 | spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_834 = 6'h27 == _T_88 | spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_835 = 6'h28 == _T_88 | spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_836 = 6'h29 == _T_88 | spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_837 = 6'h2a == _T_88 | spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_838 = 6'h2b == _T_88 | spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_839 = 6'h2c == _T_88 | spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_840 = 6'h2d == _T_88 | spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_841 = 6'h2e == _T_88 | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_842 = 6'h2f == _T_88 | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_843 = 6'h30 == _T_88 | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_844 = 6'h31 == _T_88 | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_845 = 6'h32 == _T_88 | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_846 = 6'h33 == _T_88 | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_847 = 6'h34 == _T_88 | spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_848 = 6'h35 == _T_88 | spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_849 = 6'h36 == _T_88 | spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_850 = 6'h37 == _T_88 | spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_851 = 6'h38 == _T_88 | spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_852 = 6'h39 == _T_88 | spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 471:{55,55}]
  wire  _GEN_856 = 6'h3d == _T_88 | _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 471:{55,55}]
  wire  _GEN_857 = 6'h3e == _T_88 | _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 471:{55,55}]
  wire  _GEN_858 = 6'h3f == _T_88 | _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 471:{55,55}]
  wire  _GEN_863 = _T_72 ? _GEN_798 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_864 = _T_72 ? _GEN_799 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_865 = _T_72 ? _GEN_800 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_866 = _T_72 ? _GEN_801 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_867 = _T_72 ? _GEN_802 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_868 = _T_72 ? _GEN_803 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_869 = _T_72 ? _GEN_804 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_870 = _T_72 ? _GEN_805 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_871 = _T_72 ? _GEN_806 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_872 = _T_72 ? _GEN_807 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_873 = _T_72 ? _GEN_808 : _GEN_530; // @[\\src\\main\\scala\\GameLogic.scala 470:69]
  wire  _GEN_874 = _T_72 ? _GEN_809 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_875 = _T_72 ? _GEN_810 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_876 = _T_72 ? _GEN_811 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_877 = _T_72 ? _GEN_812 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_878 = _T_72 ? _GEN_813 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_879 = _T_72 ? _GEN_814 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_880 = _T_72 ? _GEN_815 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_881 = _T_72 ? _GEN_816 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_882 = _T_72 ? _GEN_817 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_883 = _T_72 ? _GEN_818 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_884 = _T_72 ? _GEN_819 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_885 = _T_72 ? _GEN_820 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_886 = _T_72 ? _GEN_821 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_887 = _T_72 ? _GEN_822 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_888 = _T_72 ? _GEN_823 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_889 = _T_72 ? _GEN_824 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_890 = _T_72 ? _GEN_825 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_891 = _T_72 ? _GEN_826 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_892 = _T_72 ? _GEN_827 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_893 = _T_72 ? _GEN_828 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_894 = _T_72 ? _GEN_829 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_895 = _T_72 ? _GEN_830 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_896 = _T_72 ? _GEN_831 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_897 = _T_72 ? _GEN_832 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_898 = _T_72 ? _GEN_833 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_899 = _T_72 ? _GEN_834 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_900 = _T_72 ? _GEN_835 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_901 = _T_72 ? _GEN_836 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_902 = _T_72 ? _GEN_837 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_903 = _T_72 ? _GEN_838 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_904 = _T_72 ? _GEN_839 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_905 = _T_72 ? _GEN_840 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_906 = _T_72 ? _GEN_841 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_907 = _T_72 ? _GEN_842 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_908 = _T_72 ? _GEN_843 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_909 = _T_72 ? _GEN_844 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_910 = _T_72 ? _GEN_845 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_911 = _T_72 ? _GEN_846 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_912 = _T_72 ? _GEN_847 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_913 = _T_72 ? _GEN_848 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_914 = _T_72 ? _GEN_849 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_915 = _T_72 ? _GEN_850 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_916 = _T_72 ? _GEN_851 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_917 = _T_72 ? _GEN_852 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 470:69]
  wire  _GEN_921 = _T_72 ? _GEN_856 : _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 470:69]
  wire  _GEN_922 = _T_72 ? _GEN_857 : _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 470:69]
  wire  _GEN_923 = _T_72 ? _GEN_858 : _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 470:69]
  wire [7:0] _GEN_925 = _T_72 ? 8'h14 : _GEN_597; // @[\\src\\main\\scala\\GameLogic.scala 470:69 473:29]
  wire  _GEN_929 = lvlReg == 2'h3 ? _GEN_863 : spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_930 = lvlReg == 2'h3 ? _GEN_864 : spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_931 = lvlReg == 2'h3 ? _GEN_865 : spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_932 = lvlReg == 2'h3 ? _GEN_866 : spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_933 = lvlReg == 2'h3 ? _GEN_867 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_934 = lvlReg == 2'h3 ? _GEN_868 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_935 = lvlReg == 2'h3 ? _GEN_869 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_936 = lvlReg == 2'h3 ? _GEN_870 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_937 = lvlReg == 2'h3 ? _GEN_871 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_938 = lvlReg == 2'h3 ? _GEN_872 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_939 = lvlReg == 2'h3 ? _GEN_873 : _GEN_530; // @[\\src\\main\\scala\\GameLogic.scala 468:34]
  wire  _GEN_940 = lvlReg == 2'h3 ? _GEN_874 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_941 = lvlReg == 2'h3 ? _GEN_875 : spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_942 = lvlReg == 2'h3 ? _GEN_876 : spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_943 = lvlReg == 2'h3 ? _GEN_877 : spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_944 = lvlReg == 2'h3 ? _GEN_878 : spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_945 = lvlReg == 2'h3 ? _GEN_879 : spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_946 = lvlReg == 2'h3 ? _GEN_880 : spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_947 = lvlReg == 2'h3 ? _GEN_881 : spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_948 = lvlReg == 2'h3 ? _GEN_882 : spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_949 = lvlReg == 2'h3 ? _GEN_883 : spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_950 = lvlReg == 2'h3 ? _GEN_884 : spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_951 = lvlReg == 2'h3 ? _GEN_885 : spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_952 = lvlReg == 2'h3 ? _GEN_886 : spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_953 = lvlReg == 2'h3 ? _GEN_887 : spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_954 = lvlReg == 2'h3 ? _GEN_888 : spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_955 = lvlReg == 2'h3 ? _GEN_889 : spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_956 = lvlReg == 2'h3 ? _GEN_890 : spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_957 = lvlReg == 2'h3 ? _GEN_891 : spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_958 = lvlReg == 2'h3 ? _GEN_892 : spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_959 = lvlReg == 2'h3 ? _GEN_893 : spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_960 = lvlReg == 2'h3 ? _GEN_894 : spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_961 = lvlReg == 2'h3 ? _GEN_895 : spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_962 = lvlReg == 2'h3 ? _GEN_896 : spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_963 = lvlReg == 2'h3 ? _GEN_897 : spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_964 = lvlReg == 2'h3 ? _GEN_898 : spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_965 = lvlReg == 2'h3 ? _GEN_899 : spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_966 = lvlReg == 2'h3 ? _GEN_900 : spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_967 = lvlReg == 2'h3 ? _GEN_901 : spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_968 = lvlReg == 2'h3 ? _GEN_902 : spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_969 = lvlReg == 2'h3 ? _GEN_903 : spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_970 = lvlReg == 2'h3 ? _GEN_904 : spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_971 = lvlReg == 2'h3 ? _GEN_905 : spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_972 = lvlReg == 2'h3 ? _GEN_906 : spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_973 = lvlReg == 2'h3 ? _GEN_907 : spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_974 = lvlReg == 2'h3 ? _GEN_908 : spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_975 = lvlReg == 2'h3 ? _GEN_909 : spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_976 = lvlReg == 2'h3 ? _GEN_910 : spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_977 = lvlReg == 2'h3 ? _GEN_911 : spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_978 = lvlReg == 2'h3 ? _GEN_912 : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_979 = lvlReg == 2'h3 ? _GEN_913 : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_980 = lvlReg == 2'h3 ? _GEN_914 : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_981 = lvlReg == 2'h3 ? _GEN_915 : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_982 = lvlReg == 2'h3 ? _GEN_916 : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_983 = lvlReg == 2'h3 ? _GEN_917 : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 125:34 468:34]
  wire  _GEN_987 = lvlReg == 2'h3 ? _GEN_921 : _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 468:34]
  wire  _GEN_988 = lvlReg == 2'h3 ? _GEN_922 : _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 468:34]
  wire  _GEN_989 = lvlReg == 2'h3 ? _GEN_923 : _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 468:34]
  wire [5:0] _GEN_990 = lvlReg == 2'h3 ? _GEN_662 : nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 232:34 468:34]
  wire [7:0] _GEN_991 = lvlReg == 2'h3 ? _GEN_925 : spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 231:34 468:34]
  wire  _GEN_995 = lvlReg == 2'h2 ? _GEN_732 : _GEN_929; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_996 = lvlReg == 2'h2 ? _GEN_733 : _GEN_930; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_997 = lvlReg == 2'h2 ? _GEN_734 : _GEN_931; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_998 = lvlReg == 2'h2 ? _GEN_735 : _GEN_932; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_999 = lvlReg == 2'h2 ? _GEN_736 : _GEN_933; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1000 = lvlReg == 2'h2 ? _GEN_737 : _GEN_934; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1001 = lvlReg == 2'h2 ? _GEN_738 : _GEN_935; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1002 = lvlReg == 2'h2 ? _GEN_739 : _GEN_936; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1003 = lvlReg == 2'h2 ? _GEN_740 : _GEN_937; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1004 = lvlReg == 2'h2 ? _GEN_741 : _GEN_938; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1005 = lvlReg == 2'h2 ? _GEN_742 : _GEN_939; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1006 = lvlReg == 2'h2 ? _GEN_743 : _GEN_940; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1007 = lvlReg == 2'h2 ? _GEN_744 : _GEN_941; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1008 = lvlReg == 2'h2 ? _GEN_745 : _GEN_942; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1009 = lvlReg == 2'h2 ? _GEN_746 : _GEN_943; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1010 = lvlReg == 2'h2 ? _GEN_747 : _GEN_944; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1011 = lvlReg == 2'h2 ? _GEN_748 : _GEN_945; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1012 = lvlReg == 2'h2 ? _GEN_749 : _GEN_946; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1013 = lvlReg == 2'h2 ? _GEN_750 : _GEN_947; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1014 = lvlReg == 2'h2 ? _GEN_751 : _GEN_948; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1015 = lvlReg == 2'h2 ? _GEN_752 : _GEN_949; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1016 = lvlReg == 2'h2 ? _GEN_753 : _GEN_950; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1017 = lvlReg == 2'h2 ? _GEN_754 : _GEN_951; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1018 = lvlReg == 2'h2 ? _GEN_755 : _GEN_952; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1019 = lvlReg == 2'h2 ? _GEN_756 : _GEN_953; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1020 = lvlReg == 2'h2 ? _GEN_757 : _GEN_954; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1021 = lvlReg == 2'h2 ? _GEN_758 : _GEN_955; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1022 = lvlReg == 2'h2 ? _GEN_759 : _GEN_956; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1023 = lvlReg == 2'h2 ? _GEN_760 : _GEN_957; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1024 = lvlReg == 2'h2 ? _GEN_761 : _GEN_958; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1025 = lvlReg == 2'h2 ? _GEN_762 : _GEN_959; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1026 = lvlReg == 2'h2 ? _GEN_763 : _GEN_960; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1027 = lvlReg == 2'h2 ? _GEN_764 : _GEN_961; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1028 = lvlReg == 2'h2 ? _GEN_765 : _GEN_962; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1029 = lvlReg == 2'h2 ? _GEN_766 : _GEN_963; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1030 = lvlReg == 2'h2 ? _GEN_767 : _GEN_964; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1031 = lvlReg == 2'h2 ? _GEN_768 : _GEN_965; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1032 = lvlReg == 2'h2 ? _GEN_769 : _GEN_966; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1033 = lvlReg == 2'h2 ? _GEN_770 : _GEN_967; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1034 = lvlReg == 2'h2 ? _GEN_771 : _GEN_968; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1035 = lvlReg == 2'h2 ? _GEN_772 : _GEN_969; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1036 = lvlReg == 2'h2 ? _GEN_773 : _GEN_970; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1037 = lvlReg == 2'h2 ? _GEN_774 : _GEN_971; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1038 = lvlReg == 2'h2 ? _GEN_775 : _GEN_972; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1039 = lvlReg == 2'h2 ? _GEN_776 : _GEN_973; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1040 = lvlReg == 2'h2 ? _GEN_777 : _GEN_974; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1041 = lvlReg == 2'h2 ? _GEN_778 : _GEN_975; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1042 = lvlReg == 2'h2 ? _GEN_779 : _GEN_976; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1043 = lvlReg == 2'h2 ? _GEN_780 : _GEN_977; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1044 = lvlReg == 2'h2 ? _GEN_781 : _GEN_978; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1045 = lvlReg == 2'h2 ? _GEN_782 : _GEN_979; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1046 = lvlReg == 2'h2 ? _GEN_783 : _GEN_980; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1047 = lvlReg == 2'h2 ? _GEN_784 : _GEN_981; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1048 = lvlReg == 2'h2 ? _GEN_785 : _GEN_982; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1049 = lvlReg == 2'h2 ? _GEN_786 : _GEN_983; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1053 = lvlReg == 2'h2 ? _GEN_790 : _GEN_987; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1054 = lvlReg == 2'h2 ? _GEN_791 : _GEN_988; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1055 = lvlReg == 2'h2 ? _GEN_792 : _GEN_989; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire [5:0] _GEN_1056 = lvlReg == 2'h2 ? _GEN_662 : _GEN_990; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire [7:0] _GEN_1057 = lvlReg == 2'h2 ? _GEN_794 : _GEN_991; // @[\\src\\main\\scala\\GameLogic.scala 459:34]
  wire  _GEN_1071 = lvlReg == 2'h1 ? _GEN_611 : _GEN_1005; // @[\\src\\main\\scala\\GameLogic.scala 450:28]
  wire  _GEN_1072 = lvlReg == 2'h1 ? _GEN_612 : _GEN_1006; // @[\\src\\main\\scala\\GameLogic.scala 450:28]
  wire  _T_90 = ~isBlinking; // @[\\src\\main\\scala\\GameLogic.scala 482:12]
  wire [6:0] _obstacleWidth_T_1 = 5'h1a * 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 487:81]
  wire [5:0] _obstacleHeight_T_1 = 4'hf * 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 488:83]
  wire [6:0] _T_93 = spriteScaleTypeRegs_0 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2031 = {{4{_T_93[6]}},_T_93}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_96 = $signed(spriteXRegs_16) + $signed(_GEN_2031); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_97 = $signed(spriteXRegs_14) < $signed(_T_96); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_98 = spriteVisibleRegs_16 & $signed(spriteXRegs_16) <= 11'sh280 & _T_97; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [10:0] _T_101 = $signed(spriteXRegs_14) + 11'sh8; // @[\\src\\main\\scala\\GameLogic.scala 492:110]
  wire [5:0] _T_104 = spriteScaleTypeRegs_0 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2032 = {{4{_T_104[5]}},_T_104}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_107 = $signed(spriteYRegs_16) + $signed(_GEN_2032); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_108 = $signed(spriteYRegs_14) < $signed(_T_107); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_109 = _T_98 & $signed(spriteXRegs_16) < $signed(_T_101) & _T_108; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire [9:0] _T_112 = $signed(spriteYRegs_14) + 10'shb; // @[\\src\\main\\scala\\GameLogic.scala 493:111]
  wire  _T_114 = _T_109 & $signed(spriteYRegs_16) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire  _GEN_1124 = _T_114 | collisionDetected; // @[\\src\\main\\scala\\GameLogic.scala 494:13 495:31 238:34]
  wire [6:0] _T_117 = spriteScaleTypeRegs_1 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2033 = {{4{_T_117[6]}},_T_117}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_120 = $signed(spriteXRegs_17) + $signed(_GEN_2033); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_121 = $signed(spriteXRegs_14) < $signed(_T_120); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_122 = spriteVisibleRegs_17 & $signed(spriteXRegs_17) <= 11'sh280 & _T_121; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [5:0] _T_128 = spriteScaleTypeRegs_1 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2034 = {{4{_T_128[5]}},_T_128}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_131 = $signed(spriteYRegs_17) + $signed(_GEN_2034); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_132 = $signed(spriteYRegs_14) < $signed(_T_131); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_133 = _T_122 & $signed(spriteXRegs_17) < $signed(_T_101) & _T_132; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire  _T_138 = _T_133 & $signed(spriteYRegs_17) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire [6:0] _T_141 = spriteScaleTypeRegs_2 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2035 = {{4{_T_141[6]}},_T_141}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_144 = $signed(spriteXRegs_18) + $signed(_GEN_2035); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_145 = $signed(spriteXRegs_14) < $signed(_T_144); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_146 = spriteVisibleRegs_18 & $signed(spriteXRegs_18) <= 11'sh280 & _T_145; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [5:0] _T_152 = spriteScaleTypeRegs_2 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2036 = {{4{_T_152[5]}},_T_152}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_155 = $signed(spriteYRegs_18) + $signed(_GEN_2036); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_156 = $signed(spriteYRegs_14) < $signed(_T_155); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_157 = _T_146 & $signed(spriteXRegs_18) < $signed(_T_101) & _T_156; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire  _T_162 = _T_157 & $signed(spriteYRegs_18) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire [6:0] _T_165 = spriteScaleTypeRegs_3 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2037 = {{4{_T_165[6]}},_T_165}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_168 = $signed(spriteXRegs_19) + $signed(_GEN_2037); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_169 = $signed(spriteXRegs_14) < $signed(_T_168); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_170 = spriteVisibleRegs_19 & $signed(spriteXRegs_19) <= 11'sh280 & _T_169; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [5:0] _T_176 = spriteScaleTypeRegs_3 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2038 = {{4{_T_176[5]}},_T_176}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_179 = $signed(spriteYRegs_19) + $signed(_GEN_2038); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_180 = $signed(spriteYRegs_14) < $signed(_T_179); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_181 = _T_170 & $signed(spriteXRegs_19) < $signed(_T_101) & _T_180; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire  _T_186 = _T_181 & $signed(spriteYRegs_19) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire [6:0] _T_189 = spriteScaleTypeRegs_4 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2039 = {{4{_T_189[6]}},_T_189}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_192 = $signed(spriteXRegs_20) + $signed(_GEN_2039); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_193 = $signed(spriteXRegs_14) < $signed(_T_192); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_194 = spriteVisibleRegs_20 & $signed(spriteXRegs_20) <= 11'sh280 & _T_193; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [5:0] _T_200 = spriteScaleTypeRegs_4 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2040 = {{4{_T_200[5]}},_T_200}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_203 = $signed(spriteYRegs_20) + $signed(_GEN_2040); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_204 = $signed(spriteYRegs_14) < $signed(_T_203); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_205 = _T_194 & $signed(spriteXRegs_20) < $signed(_T_101) & _T_204; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire  _T_210 = _T_205 & $signed(spriteYRegs_20) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire [6:0] _T_213 = spriteScaleTypeRegs_5 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2041 = {{4{_T_213[6]}},_T_213}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_216 = $signed(spriteXRegs_21) + $signed(_GEN_2041); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_217 = $signed(spriteXRegs_14) < $signed(_T_216); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_218 = spriteVisibleRegs_21 & $signed(spriteXRegs_21) <= 11'sh280 & _T_217; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [5:0] _T_224 = spriteScaleTypeRegs_5 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2042 = {{4{_T_224[5]}},_T_224}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_227 = $signed(spriteYRegs_21) + $signed(_GEN_2042); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_228 = $signed(spriteYRegs_14) < $signed(_T_227); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_229 = _T_218 & $signed(spriteXRegs_21) < $signed(_T_101) & _T_228; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire  _T_234 = _T_229 & $signed(spriteYRegs_21) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire [6:0] _T_237 = spriteScaleTypeRegs_6 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2043 = {{4{_T_237[6]}},_T_237}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_240 = $signed(spriteXRegs_22) + $signed(_GEN_2043); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_241 = $signed(spriteXRegs_14) < $signed(_T_240); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_242 = spriteVisibleRegs_22 & $signed(spriteXRegs_22) <= 11'sh280 & _T_241; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [5:0] _T_248 = spriteScaleTypeRegs_6 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2044 = {{4{_T_248[5]}},_T_248}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_251 = $signed(spriteYRegs_22) + $signed(_GEN_2044); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_252 = $signed(spriteYRegs_14) < $signed(_T_251); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_253 = _T_242 & $signed(spriteXRegs_22) < $signed(_T_101) & _T_252; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire  _T_258 = _T_253 & $signed(spriteYRegs_22) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire [6:0] _T_261 = spriteScaleTypeRegs_7 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2045 = {{4{_T_261[6]}},_T_261}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_264 = $signed(spriteXRegs_23) + $signed(_GEN_2045); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_265 = $signed(spriteXRegs_14) < $signed(_T_264); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_266 = spriteVisibleRegs_23 & $signed(spriteXRegs_23) <= 11'sh280 & _T_265; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [5:0] _T_272 = spriteScaleTypeRegs_7 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2046 = {{4{_T_272[5]}},_T_272}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_275 = $signed(spriteYRegs_23) + $signed(_GEN_2046); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_276 = $signed(spriteYRegs_14) < $signed(_T_275); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_277 = _T_266 & $signed(spriteXRegs_23) < $signed(_T_101) & _T_276; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire  _T_282 = _T_277 & $signed(spriteYRegs_23) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire [6:0] _T_285 = spriteScaleTypeRegs_8 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2047 = {{4{_T_285[6]}},_T_285}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_288 = $signed(spriteXRegs_24) + $signed(_GEN_2047); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_289 = $signed(spriteXRegs_14) < $signed(_T_288); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_290 = spriteVisibleRegs_24 & $signed(spriteXRegs_24) <= 11'sh280 & _T_289; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [5:0] _T_296 = spriteScaleTypeRegs_8 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2048 = {{4{_T_296[5]}},_T_296}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_299 = $signed(spriteYRegs_24) + $signed(_GEN_2048); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_300 = $signed(spriteYRegs_14) < $signed(_T_299); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_301 = _T_290 & $signed(spriteXRegs_24) < $signed(_T_101) & _T_300; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire  _T_306 = _T_301 & $signed(spriteYRegs_24) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire [6:0] _T_309 = spriteScaleTypeRegs_9 ? _obstacleWidth_T_1 : 7'h1a; // @[\\src\\main\\scala\\GameLogic.scala 492:65]
  wire [10:0] _GEN_2049 = {{4{_T_309[6]}},_T_309}; // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire [10:0] _T_312 = $signed(spriteXRegs_25) + $signed(_GEN_2049); // @[\\src\\main\\scala\\GameLogic.scala 492:49]
  wire  _T_313 = $signed(spriteXRegs_14) < $signed(_T_312); // @[\\src\\main\\scala\\GameLogic.scala 492:32]
  wire  _T_314 = spriteVisibleRegs_25 & $signed(spriteXRegs_25) <= 11'sh280 & _T_313; // @[\\src\\main\\scala\\GameLogic.scala 491:63]
  wire [5:0] _T_320 = spriteScaleTypeRegs_9 ? _obstacleHeight_T_1 : 6'hf; // @[\\src\\main\\scala\\GameLogic.scala 493:66]
  wire [9:0] _GEN_2050 = {{4{_T_320[5]}},_T_320}; // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire [9:0] _T_323 = $signed(spriteYRegs_25) + $signed(_GEN_2050); // @[\\src\\main\\scala\\GameLogic.scala 493:49]
  wire  _T_324 = $signed(spriteYRegs_14) < $signed(_T_323); // @[\\src\\main\\scala\\GameLogic.scala 493:32]
  wire  _T_325 = _T_314 & $signed(spriteXRegs_25) < $signed(_T_101) & _T_324; // @[\\src\\main\\scala\\GameLogic.scala 492:117]
  wire  _T_330 = _T_325 & $signed(spriteYRegs_25) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 493:74]
  wire  _GEN_1133 = _T_330 | (_T_306 | (_T_282 | (_T_258 | (_T_234 | (_T_210 | (_T_186 | (_T_162 | (_T_138 | _GEN_1124))
    )))))); // @[\\src\\main\\scala\\GameLogic.scala 494:13 495:31]
  wire  _GEN_1134 = ~isBlinking ? _GEN_1133 : collisionDetected; // @[\\src\\main\\scala\\GameLogic.scala 482:25 238:34]
  wire [6:0] _obstacleWidth_T_21 = 5'h1d * 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 505:81]
  wire [6:0] _T_332 = spriteScaleTypeRegs_0 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2051 = {{4{_T_332[6]}},_T_332}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_335 = $signed(spriteXRegs_26) + $signed(_GEN_2051); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_336 = $signed(spriteXRegs_14) < $signed(_T_335); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_337 = spriteVisibleRegs_26 & _T_336; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_346 = $signed(spriteYRegs_26) + $signed(_GEN_2032); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_347 = $signed(spriteYRegs_14) < $signed(_T_346); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_348 = _T_337 & $signed(spriteXRegs_26) < $signed(_T_101) & _T_347; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_353 = _T_348 & $signed(spriteYRegs_26) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire [6:0] _T_354 = spriteScaleTypeRegs_1 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2053 = {{4{_T_354[6]}},_T_354}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_357 = $signed(spriteXRegs_27) + $signed(_GEN_2053); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_358 = $signed(spriteXRegs_14) < $signed(_T_357); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_359 = spriteVisibleRegs_27 & _T_358; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_368 = $signed(spriteYRegs_27) + $signed(_GEN_2034); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_369 = $signed(spriteYRegs_14) < $signed(_T_368); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_370 = _T_359 & $signed(spriteXRegs_27) < $signed(_T_101) & _T_369; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_375 = _T_370 & $signed(spriteYRegs_27) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire [6:0] _T_376 = spriteScaleTypeRegs_2 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2055 = {{4{_T_376[6]}},_T_376}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_379 = $signed(spriteXRegs_28) + $signed(_GEN_2055); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_380 = $signed(spriteXRegs_14) < $signed(_T_379); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_381 = spriteVisibleRegs_28 & _T_380; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_390 = $signed(spriteYRegs_28) + $signed(_GEN_2036); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_391 = $signed(spriteYRegs_14) < $signed(_T_390); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_392 = _T_381 & $signed(spriteXRegs_28) < $signed(_T_101) & _T_391; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_397 = _T_392 & $signed(spriteYRegs_28) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire [6:0] _T_398 = spriteScaleTypeRegs_3 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2057 = {{4{_T_398[6]}},_T_398}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_401 = $signed(spriteXRegs_29) + $signed(_GEN_2057); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_402 = $signed(spriteXRegs_14) < $signed(_T_401); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_403 = spriteVisibleRegs_29 & _T_402; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_412 = $signed(spriteYRegs_29) + $signed(_GEN_2038); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_413 = $signed(spriteYRegs_14) < $signed(_T_412); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_414 = _T_403 & $signed(spriteXRegs_29) < $signed(_T_101) & _T_413; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_419 = _T_414 & $signed(spriteYRegs_29) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire [6:0] _T_420 = spriteScaleTypeRegs_4 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2059 = {{4{_T_420[6]}},_T_420}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_423 = $signed(spriteXRegs_30) + $signed(_GEN_2059); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_424 = $signed(spriteXRegs_14) < $signed(_T_423); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_425 = spriteVisibleRegs_30 & _T_424; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_434 = $signed(spriteYRegs_30) + $signed(_GEN_2040); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_435 = $signed(spriteYRegs_14) < $signed(_T_434); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_436 = _T_425 & $signed(spriteXRegs_30) < $signed(_T_101) & _T_435; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_441 = _T_436 & $signed(spriteYRegs_30) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire [6:0] _T_442 = spriteScaleTypeRegs_5 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2061 = {{4{_T_442[6]}},_T_442}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_445 = $signed(spriteXRegs_31) + $signed(_GEN_2061); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_446 = $signed(spriteXRegs_14) < $signed(_T_445); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_447 = spriteVisibleRegs_31 & _T_446; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_456 = $signed(spriteYRegs_31) + $signed(_GEN_2042); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_457 = $signed(spriteYRegs_14) < $signed(_T_456); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_458 = _T_447 & $signed(spriteXRegs_31) < $signed(_T_101) & _T_457; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_463 = _T_458 & $signed(spriteYRegs_31) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire [6:0] _T_464 = spriteScaleTypeRegs_6 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2063 = {{4{_T_464[6]}},_T_464}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_467 = $signed(spriteXRegs_32) + $signed(_GEN_2063); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_468 = $signed(spriteXRegs_14) < $signed(_T_467); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_469 = spriteVisibleRegs_32 & _T_468; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_478 = $signed(spriteYRegs_32) + $signed(_GEN_2044); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_479 = $signed(spriteYRegs_14) < $signed(_T_478); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_480 = _T_469 & $signed(spriteXRegs_32) < $signed(_T_101) & _T_479; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_485 = _T_480 & $signed(spriteYRegs_32) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire [6:0] _T_486 = spriteScaleTypeRegs_7 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2065 = {{4{_T_486[6]}},_T_486}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_489 = $signed(spriteXRegs_33) + $signed(_GEN_2065); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_490 = $signed(spriteXRegs_14) < $signed(_T_489); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_491 = spriteVisibleRegs_33 & _T_490; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_500 = $signed(spriteYRegs_33) + $signed(_GEN_2046); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_501 = $signed(spriteYRegs_14) < $signed(_T_500); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_502 = _T_491 & $signed(spriteXRegs_33) < $signed(_T_101) & _T_501; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_507 = _T_502 & $signed(spriteYRegs_33) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire [6:0] _T_508 = spriteScaleTypeRegs_8 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2067 = {{4{_T_508[6]}},_T_508}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_511 = $signed(spriteXRegs_34) + $signed(_GEN_2067); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_512 = $signed(spriteXRegs_14) < $signed(_T_511); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_513 = spriteVisibleRegs_34 & _T_512; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_522 = $signed(spriteYRegs_34) + $signed(_GEN_2048); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_523 = $signed(spriteYRegs_14) < $signed(_T_522); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_524 = _T_513 & $signed(spriteXRegs_34) < $signed(_T_101) & _T_523; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_529 = _T_524 & $signed(spriteYRegs_34) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire [6:0] _T_530 = spriteScaleTypeRegs_9 ? _obstacleWidth_T_21 : 7'h1d; // @[\\src\\main\\scala\\GameLogic.scala 510:65]
  wire [10:0] _GEN_2069 = {{4{_T_530[6]}},_T_530}; // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire [10:0] _T_533 = $signed(spriteXRegs_35) + $signed(_GEN_2069); // @[\\src\\main\\scala\\GameLogic.scala 510:49]
  wire  _T_534 = $signed(spriteXRegs_14) < $signed(_T_533); // @[\\src\\main\\scala\\GameLogic.scala 510:32]
  wire  _T_535 = spriteVisibleRegs_35 & _T_534; // @[\\src\\main\\scala\\GameLogic.scala 509:34]
  wire [9:0] _T_544 = $signed(spriteYRegs_35) + $signed(_GEN_2050); // @[\\src\\main\\scala\\GameLogic.scala 511:49]
  wire  _T_545 = $signed(spriteYRegs_14) < $signed(_T_544); // @[\\src\\main\\scala\\GameLogic.scala 511:32]
  wire  _T_546 = _T_535 & $signed(spriteXRegs_35) < $signed(_T_101) & _T_545; // @[\\src\\main\\scala\\GameLogic.scala 510:117]
  wire  _T_551 = _T_546 & $signed(spriteYRegs_35) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 511:74]
  wire  _GEN_1144 = _T_551 | (_T_529 | (_T_507 | (_T_485 | (_T_463 | (_T_441 | (_T_419 | (_T_397 | (_T_375 | (_T_353 |
    _GEN_1134))))))))); // @[\\src\\main\\scala\\GameLogic.scala 512:13 513:31]
  wire  _GEN_1145 = _T_90 ? _GEN_1144 : _GEN_1134; // @[\\src\\main\\scala\\GameLogic.scala 500:25]
  wire [7:0] _obstacleWidth_T_41 = 6'h20 * 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 523:81]
  wire [7:0] _T_553 = spriteScaleTypeRegs_0 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2071 = {{3{_T_553[7]}},_T_553}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_556 = $signed(spriteXRegs_36) + $signed(_GEN_2071); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_557 = $signed(spriteXRegs_14) < $signed(_T_556); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_558 = spriteVisibleRegs_36 & _T_557; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_567 = $signed(spriteYRegs_36) + $signed(_GEN_2032); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_568 = $signed(spriteYRegs_14) < $signed(_T_567); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_569 = _T_558 & $signed(spriteXRegs_36) < $signed(_T_101) & _T_568; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_574 = _T_569 & $signed(spriteYRegs_36) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire [7:0] _T_575 = spriteScaleTypeRegs_1 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2073 = {{3{_T_575[7]}},_T_575}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_578 = $signed(spriteXRegs_37) + $signed(_GEN_2073); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_579 = $signed(spriteXRegs_14) < $signed(_T_578); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_580 = spriteVisibleRegs_37 & _T_579; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_589 = $signed(spriteYRegs_37) + $signed(_GEN_2034); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_590 = $signed(spriteYRegs_14) < $signed(_T_589); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_591 = _T_580 & $signed(spriteXRegs_37) < $signed(_T_101) & _T_590; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_596 = _T_591 & $signed(spriteYRegs_37) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire [7:0] _T_597 = spriteScaleTypeRegs_2 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2075 = {{3{_T_597[7]}},_T_597}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_600 = $signed(spriteXRegs_38) + $signed(_GEN_2075); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_601 = $signed(spriteXRegs_14) < $signed(_T_600); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_602 = spriteVisibleRegs_38 & _T_601; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_611 = $signed(spriteYRegs_38) + $signed(_GEN_2036); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_612 = $signed(spriteYRegs_14) < $signed(_T_611); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_613 = _T_602 & $signed(spriteXRegs_38) < $signed(_T_101) & _T_612; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_618 = _T_613 & $signed(spriteYRegs_38) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire [7:0] _T_619 = spriteScaleTypeRegs_3 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2077 = {{3{_T_619[7]}},_T_619}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_622 = $signed(spriteXRegs_39) + $signed(_GEN_2077); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_623 = $signed(spriteXRegs_14) < $signed(_T_622); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_624 = spriteVisibleRegs_39 & _T_623; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_633 = $signed(spriteYRegs_39) + $signed(_GEN_2038); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_634 = $signed(spriteYRegs_14) < $signed(_T_633); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_635 = _T_624 & $signed(spriteXRegs_39) < $signed(_T_101) & _T_634; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_640 = _T_635 & $signed(spriteYRegs_39) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire [7:0] _T_641 = spriteScaleTypeRegs_4 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2079 = {{3{_T_641[7]}},_T_641}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_644 = $signed(spriteXRegs_40) + $signed(_GEN_2079); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_645 = $signed(spriteXRegs_14) < $signed(_T_644); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_646 = spriteVisibleRegs_40 & _T_645; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_655 = $signed(spriteYRegs_40) + $signed(_GEN_2040); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_656 = $signed(spriteYRegs_14) < $signed(_T_655); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_657 = _T_646 & $signed(spriteXRegs_40) < $signed(_T_101) & _T_656; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_662 = _T_657 & $signed(spriteYRegs_40) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire [7:0] _T_663 = spriteScaleTypeRegs_5 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2081 = {{3{_T_663[7]}},_T_663}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_666 = $signed(spriteXRegs_41) + $signed(_GEN_2081); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_667 = $signed(spriteXRegs_14) < $signed(_T_666); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_668 = spriteVisibleRegs_41 & _T_667; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_677 = $signed(spriteYRegs_41) + $signed(_GEN_2042); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_678 = $signed(spriteYRegs_14) < $signed(_T_677); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_679 = _T_668 & $signed(spriteXRegs_41) < $signed(_T_101) & _T_678; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_684 = _T_679 & $signed(spriteYRegs_41) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire [7:0] _T_685 = spriteScaleTypeRegs_6 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2083 = {{3{_T_685[7]}},_T_685}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_688 = $signed(spriteXRegs_42) + $signed(_GEN_2083); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_689 = $signed(spriteXRegs_14) < $signed(_T_688); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_690 = spriteVisibleRegs_42 & _T_689; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_699 = $signed(spriteYRegs_42) + $signed(_GEN_2044); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_700 = $signed(spriteYRegs_14) < $signed(_T_699); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_701 = _T_690 & $signed(spriteXRegs_42) < $signed(_T_101) & _T_700; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_706 = _T_701 & $signed(spriteYRegs_42) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire [7:0] _T_707 = spriteScaleTypeRegs_7 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2085 = {{3{_T_707[7]}},_T_707}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_710 = $signed(spriteXRegs_43) + $signed(_GEN_2085); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_711 = $signed(spriteXRegs_14) < $signed(_T_710); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_712 = spriteVisibleRegs_43 & _T_711; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_721 = $signed(spriteYRegs_43) + $signed(_GEN_2046); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_722 = $signed(spriteYRegs_14) < $signed(_T_721); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_723 = _T_712 & $signed(spriteXRegs_43) < $signed(_T_101) & _T_722; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_728 = _T_723 & $signed(spriteYRegs_43) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire [7:0] _T_729 = spriteScaleTypeRegs_8 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2087 = {{3{_T_729[7]}},_T_729}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_732 = $signed(spriteXRegs_44) + $signed(_GEN_2087); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_733 = $signed(spriteXRegs_14) < $signed(_T_732); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_734 = spriteVisibleRegs_44 & _T_733; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_743 = $signed(spriteYRegs_44) + $signed(_GEN_2048); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_744 = $signed(spriteYRegs_14) < $signed(_T_743); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_745 = _T_734 & $signed(spriteXRegs_44) < $signed(_T_101) & _T_744; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_750 = _T_745 & $signed(spriteYRegs_44) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire [7:0] _T_751 = spriteScaleTypeRegs_9 ? _obstacleWidth_T_41 : 8'h20; // @[\\src\\main\\scala\\GameLogic.scala 527:65]
  wire [10:0] _GEN_2089 = {{3{_T_751[7]}},_T_751}; // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire [10:0] _T_754 = $signed(spriteXRegs_45) + $signed(_GEN_2089); // @[\\src\\main\\scala\\GameLogic.scala 527:49]
  wire  _T_755 = $signed(spriteXRegs_14) < $signed(_T_754); // @[\\src\\main\\scala\\GameLogic.scala 527:32]
  wire  _T_756 = spriteVisibleRegs_45 & _T_755; // @[\\src\\main\\scala\\GameLogic.scala 526:34]
  wire [9:0] _T_765 = $signed(spriteYRegs_45) + $signed(_GEN_2050); // @[\\src\\main\\scala\\GameLogic.scala 528:49]
  wire  _T_766 = $signed(spriteYRegs_14) < $signed(_T_765); // @[\\src\\main\\scala\\GameLogic.scala 528:32]
  wire  _T_767 = _T_756 & $signed(spriteXRegs_45) < $signed(_T_101) & _T_766; // @[\\src\\main\\scala\\GameLogic.scala 527:117]
  wire  _T_772 = _T_767 & $signed(spriteYRegs_45) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 528:74]
  wire  _GEN_1155 = _T_772 | (_T_750 | (_T_728 | (_T_706 | (_T_684 | (_T_662 | (_T_640 | (_T_618 | (_T_596 | (_T_574 |
    _GEN_1145))))))))); // @[\\src\\main\\scala\\GameLogic.scala 529:13 530:31]
  wire  _GEN_1156 = _T_90 ? _GEN_1155 : _GEN_1145; // @[\\src\\main\\scala\\GameLogic.scala 518:25]
  wire [10:0] _T_775 = $signed(spriteXRegs_13) + 11'sh16; // @[\\src\\main\\scala\\GameLogic.scala 538:46]
  wire  _T_776 = $signed(spriteXRegs_14) < $signed(_T_775); // @[\\src\\main\\scala\\GameLogic.scala 538:28]
  wire  _T_777 = spriteVisibleRegs_13 & _T_776; // @[\\src\\main\\scala\\GameLogic.scala 537:31]
  wire [9:0] _T_785 = $signed(spriteYRegs_13) + 10'sh16; // @[\\src\\main\\scala\\GameLogic.scala 539:46]
  wire  _T_786 = $signed(spriteYRegs_14) < $signed(_T_785); // @[\\src\\main\\scala\\GameLogic.scala 539:28]
  wire  _T_787 = _T_777 & $signed(spriteXRegs_13) < $signed(_T_101) & _T_786; // @[\\src\\main\\scala\\GameLogic.scala 538:99]
  wire  _T_792 = _T_787 & $signed(spriteYRegs_13) < $signed(_T_112); // @[\\src\\main\\scala\\GameLogic.scala 539:54]
  wire [2:0] _livesReg_T_1 = livesReg + 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 543:32]
  wire [2:0] _GEN_1157 = livesReg < 3'h3 ? _livesReg_T_1 : livesReg; // @[\\src\\main\\scala\\GameLogic.scala 542:30 543:20 222:25]
  wire [2:0] _GEN_1159 = _T_792 ? _GEN_1157 : livesReg; // @[\\src\\main\\scala\\GameLogic.scala 222:25 540:9]
  wire  _GEN_1160 = collisionDetected & _T_90 | isBlinking; // @[\\src\\main\\scala\\GameLogic.scala 548:46 549:20 241:27]
  wire [7:0] _GEN_1161 = collisionDetected & _T_90 ? 8'h0 : blinkCounter; // @[\\src\\main\\scala\\GameLogic.scala 548:46 550:22 239:29]
  wire [1:0] _GEN_1162 = collisionDetected & _T_90 ? 2'h0 : blinkTimes; // @[\\src\\main\\scala\\GameLogic.scala 548:46 551:20 240:27]
  wire  _GEN_1163 = blinkCounter < 8'h14 | _GEN_1072; // @[\\src\\main\\scala\\GameLogic.scala 559:41 560:33]
  wire  _GEN_1164 = blinkCounter < 8'ha ? 1'h0 : _GEN_1163; // @[\\src\\main\\scala\\GameLogic.scala 557:35 558:33]
  wire [7:0] _blinkCounter_T_1 = blinkCounter + 8'h1; // @[\\src\\main\\scala\\GameLogic.scala 562:38]
  wire [1:0] _blinkTimes_T_1 = blinkTimes + 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 565:36]
  wire [7:0] _GEN_1165 = blinkCounter == 8'h14 ? 8'h0 : _blinkCounter_T_1; // @[\\src\\main\\scala\\GameLogic.scala 562:22 563:37 564:24]
  wire [1:0] _GEN_1166 = blinkCounter == 8'h14 ? _blinkTimes_T_1 : _GEN_1162; // @[\\src\\main\\scala\\GameLogic.scala 563:37 565:22]
  wire [2:0] _livesReg_T_3 = livesReg - 3'h1; // @[\\src\\main\\scala\\GameLogic.scala 574:34]
  wire [2:0] _GEN_1167 = livesReg <= 3'h1 ? 3'h0 : _livesReg_T_3; // @[\\src\\main\\scala\\GameLogic.scala 570:33 571:22 574:22]
  wire [2:0] _GEN_1168 = livesReg <= 3'h1 ? 3'h6 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 570:33 572:22 113:25]
  wire  _GEN_1169 = blinkTimes == 2'h3 ? 1'h0 : _GEN_1160; // @[\\src\\main\\scala\\GameLogic.scala 567:34 568:22]
  wire  _GEN_1170 = blinkTimes == 2'h3 | _GEN_1164; // @[\\src\\main\\scala\\GameLogic.scala 567:34 569:33]
  wire [2:0] _GEN_1171 = blinkTimes == 2'h3 ? _GEN_1167 : _GEN_1159; // @[\\src\\main\\scala\\GameLogic.scala 567:34]
  wire [2:0] _GEN_1172 = blinkTimes == 2'h3 ? _GEN_1168 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 113:25 567:34]
  wire  _GEN_1173 = blinkTimes == 2'h3 ? 1'h0 : _GEN_1156; // @[\\src\\main\\scala\\GameLogic.scala 567:34 576:29]
  wire [2:0] _GEN_1179 = isBlinking ? _GEN_1172 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 555:24 113:25]
  reg [10:0] spriteXRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 595:35]
  reg [9:0] spriteYRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 596:35]
  reg [10:0] spriteXRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 597:35]
  reg [9:0] spriteYRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 598:35]
  reg [10:0] spriteXRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 599:35]
  reg [9:0] spriteYRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 600:35]
  wire [9:0] _starCnt_T_1 = starCnt + 10'h1; // @[\\src\\main\\scala\\GameLogic.scala 607:28]
  wire [10:0] _spriteXRegs_58_T_5 = $signed(spriteXRegs_58) + 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 615:44]
  wire [10:0] _spriteXRegs_59_T_5 = $signed(spriteXRegs_59) + 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 616:44]
  wire [10:0] _spriteXRegs_60_T_5 = $signed(spriteXRegs_60) + 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 617:44]
  wire [9:0] _spriteYRegs_58_T_5 = $signed(spriteYRegs_58) + 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 618:44]
  wire [9:0] _spriteYRegs_59_T_5 = $signed(spriteYRegs_59) + 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 619:44]
  wire [9:0] _spriteYRegs_60_T_5 = $signed(spriteYRegs_60) + 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 620:44]
  reg [10:0] spriteXRegs_58_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 623:35]
  reg [9:0] spriteYRegs_58_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 624:35]
  reg [10:0] spriteXRegs_59_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 625:35]
  reg [9:0] spriteYRegs_59_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 626:35]
  reg [10:0] spriteXRegs_60_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 627:35]
  reg [9:0] spriteYRegs_60_REG_1; // @[\\src\\main\\scala\\GameLogic.scala 628:35]
  reg [10:0] spriteXRegs_58_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 651:35]
  reg [9:0] spriteYRegs_58_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 652:35]
  reg [10:0] spriteXRegs_59_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 653:35]
  reg [9:0] spriteYRegs_59_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 654:35]
  reg [10:0] spriteXRegs_60_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 655:35]
  reg [9:0] spriteYRegs_60_REG_2; // @[\\src\\main\\scala\\GameLogic.scala 656:35]
  wire [9:0] _GEN_1182 = starCnt == 10'h168 ? 10'h0 : _starCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 678:37 679:17 681:17]
  wire  _GEN_1183 = starCnt == 10'h12c ? 1'h0 : sprite58ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 664:37 665:35 168:42]
  wire  _GEN_1184 = starCnt == 10'h12c ? 1'h0 : sprite59ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 664:37 666:35 170:42]
  wire  _GEN_1185 = starCnt == 10'h12c ? 1'h0 : sprite60ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 664:37 667:35 172:42]
  wire  _GEN_1186 = starCnt == 10'h12c ? 1'h0 : sprite58ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 664:37 668:33 169:40]
  wire  _GEN_1187 = starCnt == 10'h12c ? 1'h0 : sprite59ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 664:37 669:33 171:40]
  wire  _GEN_1188 = starCnt == 10'h12c ? 1'h0 : sprite60ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 664:37 670:33 173:40]
  wire [10:0] _GEN_1189 = starCnt == 10'h12c ? $signed(_spriteXRegs_58_T_5) : $signed(_GEN_102); // @[\\src\\main\\scala\\GameLogic.scala 664:37 671:25]
  wire [10:0] _GEN_1190 = starCnt == 10'h12c ? $signed(_spriteXRegs_59_T_5) : $signed(_GEN_104); // @[\\src\\main\\scala\\GameLogic.scala 664:37 672:25]
  wire [10:0] _GEN_1191 = starCnt == 10'h12c ? $signed(_spriteXRegs_60_T_5) : $signed(_GEN_106); // @[\\src\\main\\scala\\GameLogic.scala 664:37 673:25]
  wire [9:0] _GEN_1192 = starCnt == 10'h12c ? $signed(_spriteYRegs_58_T_5) : $signed(_GEN_103); // @[\\src\\main\\scala\\GameLogic.scala 664:37 674:25]
  wire [9:0] _GEN_1193 = starCnt == 10'h12c ? $signed(_spriteYRegs_59_T_5) : $signed(_GEN_105); // @[\\src\\main\\scala\\GameLogic.scala 664:37 675:25]
  wire [9:0] _GEN_1194 = starCnt == 10'h12c ? $signed(_spriteYRegs_60_T_5) : $signed(_GEN_107); // @[\\src\\main\\scala\\GameLogic.scala 664:37 676:25]
  wire [9:0] _GEN_1195 = starCnt == 10'h12c ? _starCnt_T_1 : _GEN_1182; // @[\\src\\main\\scala\\GameLogic.scala 664:37 677:17]
  wire [10:0] _GEN_1196 = starCnt == 10'hf0 ? $signed(spriteXRegs_58_REG_2) : $signed(_GEN_1189); // @[\\src\\main\\scala\\GameLogic.scala 650:37 651:25]
  wire [9:0] _GEN_1197 = starCnt == 10'hf0 ? $signed(spriteYRegs_58_REG_2) : $signed(_GEN_1192); // @[\\src\\main\\scala\\GameLogic.scala 650:37 652:25]
  wire [10:0] _GEN_1198 = starCnt == 10'hf0 ? $signed(spriteXRegs_59_REG_2) : $signed(_GEN_1190); // @[\\src\\main\\scala\\GameLogic.scala 650:37 653:25]
  wire [9:0] _GEN_1199 = starCnt == 10'hf0 ? $signed(spriteYRegs_59_REG_2) : $signed(_GEN_1193); // @[\\src\\main\\scala\\GameLogic.scala 650:37 654:25]
  wire [10:0] _GEN_1200 = starCnt == 10'hf0 ? $signed(spriteXRegs_60_REG_2) : $signed(_GEN_1191); // @[\\src\\main\\scala\\GameLogic.scala 650:37 655:25]
  wire [9:0] _GEN_1201 = starCnt == 10'hf0 ? $signed(spriteYRegs_60_REG_2) : $signed(_GEN_1194); // @[\\src\\main\\scala\\GameLogic.scala 650:37 656:25]
  wire  _GEN_1202 = starCnt == 10'hf0 | _GEN_1183; // @[\\src\\main\\scala\\GameLogic.scala 650:37 657:35]
  wire  _GEN_1203 = starCnt == 10'hf0 | _GEN_1184; // @[\\src\\main\\scala\\GameLogic.scala 650:37 658:35]
  wire  _GEN_1204 = starCnt == 10'hf0 | _GEN_1185; // @[\\src\\main\\scala\\GameLogic.scala 650:37 659:35]
  wire  _GEN_1205 = starCnt == 10'hf0 | _GEN_1186; // @[\\src\\main\\scala\\GameLogic.scala 650:37 660:33]
  wire  _GEN_1206 = starCnt == 10'hf0 | _GEN_1187; // @[\\src\\main\\scala\\GameLogic.scala 650:37 661:33]
  wire  _GEN_1207 = starCnt == 10'hf0 | _GEN_1188; // @[\\src\\main\\scala\\GameLogic.scala 650:37 662:33]
  wire [9:0] _GEN_1208 = starCnt == 10'hf0 ? _starCnt_T_1 : _GEN_1195; // @[\\src\\main\\scala\\GameLogic.scala 650:37 663:17]
  wire  _GEN_1209 = starCnt == 10'hb4 ? 1'h0 : _GEN_1202; // @[\\src\\main\\scala\\GameLogic.scala 636:37 637:35]
  wire  _GEN_1210 = starCnt == 10'hb4 ? 1'h0 : _GEN_1203; // @[\\src\\main\\scala\\GameLogic.scala 636:37 638:35]
  wire  _GEN_1211 = starCnt == 10'hb4 ? 1'h0 : _GEN_1204; // @[\\src\\main\\scala\\GameLogic.scala 636:37 639:35]
  wire  _GEN_1212 = starCnt == 10'hb4 ? 1'h0 : _GEN_1205; // @[\\src\\main\\scala\\GameLogic.scala 636:37 640:33]
  wire  _GEN_1213 = starCnt == 10'hb4 ? 1'h0 : _GEN_1206; // @[\\src\\main\\scala\\GameLogic.scala 636:37 641:33]
  wire  _GEN_1214 = starCnt == 10'hb4 ? 1'h0 : _GEN_1207; // @[\\src\\main\\scala\\GameLogic.scala 636:37 642:33]
  wire [10:0] _GEN_1215 = starCnt == 10'hb4 ? $signed(_spriteXRegs_58_T_5) : $signed(_GEN_1196); // @[\\src\\main\\scala\\GameLogic.scala 636:37 643:25]
  wire [10:0] _GEN_1216 = starCnt == 10'hb4 ? $signed(_spriteXRegs_59_T_5) : $signed(_GEN_1198); // @[\\src\\main\\scala\\GameLogic.scala 636:37 644:25]
  wire [10:0] _GEN_1217 = starCnt == 10'hb4 ? $signed(_spriteXRegs_60_T_5) : $signed(_GEN_1200); // @[\\src\\main\\scala\\GameLogic.scala 636:37 645:25]
  wire [9:0] _GEN_1218 = starCnt == 10'hb4 ? $signed(_spriteYRegs_58_T_5) : $signed(_GEN_1197); // @[\\src\\main\\scala\\GameLogic.scala 636:37 646:25]
  wire [9:0] _GEN_1219 = starCnt == 10'hb4 ? $signed(_spriteYRegs_59_T_5) : $signed(_GEN_1199); // @[\\src\\main\\scala\\GameLogic.scala 636:37 647:25]
  wire [9:0] _GEN_1220 = starCnt == 10'hb4 ? $signed(_spriteYRegs_60_T_5) : $signed(_GEN_1201); // @[\\src\\main\\scala\\GameLogic.scala 636:37 648:25]
  wire [9:0] _GEN_1221 = starCnt == 10'hb4 ? _starCnt_T_1 : _GEN_1208; // @[\\src\\main\\scala\\GameLogic.scala 636:37 649:17]
  wire [10:0] _GEN_1222 = starCnt == 10'h78 ? $signed(spriteXRegs_58_REG_1) : $signed(_GEN_1215); // @[\\src\\main\\scala\\GameLogic.scala 622:37 623:25]
  wire [9:0] _GEN_1223 = starCnt == 10'h78 ? $signed(spriteYRegs_58_REG_1) : $signed(_GEN_1218); // @[\\src\\main\\scala\\GameLogic.scala 622:37 624:25]
  wire [10:0] _GEN_1224 = starCnt == 10'h78 ? $signed(spriteXRegs_59_REG_1) : $signed(_GEN_1216); // @[\\src\\main\\scala\\GameLogic.scala 622:37 625:25]
  wire [9:0] _GEN_1225 = starCnt == 10'h78 ? $signed(spriteYRegs_59_REG_1) : $signed(_GEN_1219); // @[\\src\\main\\scala\\GameLogic.scala 622:37 626:25]
  wire [10:0] _GEN_1226 = starCnt == 10'h78 ? $signed(spriteXRegs_60_REG_1) : $signed(_GEN_1217); // @[\\src\\main\\scala\\GameLogic.scala 622:37 627:25]
  wire [9:0] _GEN_1227 = starCnt == 10'h78 ? $signed(spriteYRegs_60_REG_1) : $signed(_GEN_1220); // @[\\src\\main\\scala\\GameLogic.scala 622:37 628:25]
  wire  _GEN_1228 = starCnt == 10'h78 | _GEN_1209; // @[\\src\\main\\scala\\GameLogic.scala 622:37 629:35]
  wire  _GEN_1229 = starCnt == 10'h78 | _GEN_1210; // @[\\src\\main\\scala\\GameLogic.scala 622:37 630:35]
  wire  _GEN_1230 = starCnt == 10'h78 | _GEN_1211; // @[\\src\\main\\scala\\GameLogic.scala 622:37 631:35]
  wire  _GEN_1231 = starCnt == 10'h78 | _GEN_1212; // @[\\src\\main\\scala\\GameLogic.scala 622:37 632:33]
  wire  _GEN_1232 = starCnt == 10'h78 | _GEN_1213; // @[\\src\\main\\scala\\GameLogic.scala 622:37 633:33]
  wire  _GEN_1233 = starCnt == 10'h78 | _GEN_1214; // @[\\src\\main\\scala\\GameLogic.scala 622:37 634:33]
  wire [9:0] _GEN_1234 = starCnt == 10'h78 ? _starCnt_T_1 : _GEN_1221; // @[\\src\\main\\scala\\GameLogic.scala 622:37 635:17]
  wire  _GEN_1235 = starCnt == 10'h3c ? 1'h0 : _GEN_1228; // @[\\src\\main\\scala\\GameLogic.scala 608:36 609:35]
  wire  _GEN_1236 = starCnt == 10'h3c ? 1'h0 : _GEN_1229; // @[\\src\\main\\scala\\GameLogic.scala 608:36 610:35]
  wire  _GEN_1237 = starCnt == 10'h3c ? 1'h0 : _GEN_1230; // @[\\src\\main\\scala\\GameLogic.scala 608:36 611:35]
  wire  _GEN_1238 = starCnt == 10'h3c ? 1'h0 : _GEN_1231; // @[\\src\\main\\scala\\GameLogic.scala 608:36 612:33]
  wire  _GEN_1239 = starCnt == 10'h3c ? 1'h0 : _GEN_1232; // @[\\src\\main\\scala\\GameLogic.scala 608:36 613:33]
  wire  _GEN_1240 = starCnt == 10'h3c ? 1'h0 : _GEN_1233; // @[\\src\\main\\scala\\GameLogic.scala 608:36 614:33]
  wire [10:0] _GEN_1241 = starCnt == 10'h3c ? $signed(_spriteXRegs_58_T_5) : $signed(_GEN_1222); // @[\\src\\main\\scala\\GameLogic.scala 608:36 615:25]
  wire [10:0] _GEN_1242 = starCnt == 10'h3c ? $signed(_spriteXRegs_59_T_5) : $signed(_GEN_1224); // @[\\src\\main\\scala\\GameLogic.scala 608:36 616:25]
  wire [10:0] _GEN_1243 = starCnt == 10'h3c ? $signed(_spriteXRegs_60_T_5) : $signed(_GEN_1226); // @[\\src\\main\\scala\\GameLogic.scala 608:36 617:25]
  wire [9:0] _GEN_1244 = starCnt == 10'h3c ? $signed(_spriteYRegs_58_T_5) : $signed(_GEN_1223); // @[\\src\\main\\scala\\GameLogic.scala 608:36 618:25]
  wire [9:0] _GEN_1245 = starCnt == 10'h3c ? $signed(_spriteYRegs_59_T_5) : $signed(_GEN_1225); // @[\\src\\main\\scala\\GameLogic.scala 608:36 619:25]
  wire [9:0] _GEN_1246 = starCnt == 10'h3c ? $signed(_spriteYRegs_60_T_5) : $signed(_GEN_1227); // @[\\src\\main\\scala\\GameLogic.scala 608:36 620:25]
  wire [9:0] _GEN_1247 = starCnt == 10'h3c ? _starCnt_T_1 : _GEN_1234; // @[\\src\\main\\scala\\GameLogic.scala 608:36 621:17]
  wire  _GEN_1254 = starCnt == 10'h0 | _GEN_1235; // @[\\src\\main\\scala\\GameLogic.scala 594:29 601:35]
  wire  _GEN_1255 = starCnt == 10'h0 | _GEN_1236; // @[\\src\\main\\scala\\GameLogic.scala 594:29 602:35]
  wire  _GEN_1256 = starCnt == 10'h0 | _GEN_1237; // @[\\src\\main\\scala\\GameLogic.scala 594:29 603:35]
  wire  _GEN_1257 = starCnt == 10'h0 | _GEN_1238; // @[\\src\\main\\scala\\GameLogic.scala 594:29 604:33]
  wire  _GEN_1258 = starCnt == 10'h0 | _GEN_1239; // @[\\src\\main\\scala\\GameLogic.scala 594:29 605:33]
  wire  _GEN_1259 = starCnt == 10'h0 | _GEN_1240; // @[\\src\\main\\scala\\GameLogic.scala 594:29 606:33]
  wire  _T_815 = $signed(spriteYRegs_3) > 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 702:81]
  wire  _T_817 = $signed(spriteYRegs_3) < 10'sh14c; // @[\\src\\main\\scala\\GameLogic.scala 702:107]
  wire  _T_818 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c; // @[\\src\\main\\scala\\GameLogic.scala 702:89]
  wire [1:0] _GEN_1262 = io_btnC ? 2'h1 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 705:25 706:20 211:23]
  wire [2:0] _GEN_1263 = io_btnC ? 3'h3 : 3'h4; // @[\\src\\main\\scala\\GameLogic.scala 705:25 707:22 709:22]
  wire  _T_825 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817; // @[\\src\\main\\scala\\GameLogic.scala 711:95]
  wire [1:0] _GEN_1264 = io_btnC ? 2'h2 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 714:25 715:20 211:23]
  wire  _T_832 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_815 & _T_817; // @[\\src\\main\\scala\\GameLogic.scala 720:95]
  wire [1:0] _GEN_1265 = io_btnC ? 2'h3 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 723:25 724:20 211:23]
  wire  _GEN_1266 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_815 & _T_817 ? 1'h0 : 1'h1
    ; // @[\\src\\main\\scala\\GameLogic.scala 720:122 699:31 721:33]
  wire [1:0] _GEN_1268 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_815 & _T_817 ?
    _GEN_1265 : lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 720:122 211:23]
  wire [2:0] _GEN_1269 = $signed(spriteXRegs_3) > 11'sh143 & $signed(spriteXRegs_3) < 11'sh163 & _T_815 & _T_817 ?
    _GEN_1263 : 3'h4; // @[\\src\\main\\scala\\GameLogic.scala 720:122 730:20]
  wire  _GEN_1270 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 ? 1'h0 : 1'h1
    ; // @[\\src\\main\\scala\\GameLogic.scala 711:122 697:30 712:32]
  wire [1:0] _GEN_1272 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 ?
    _GEN_1264 : _GEN_1268; // @[\\src\\main\\scala\\GameLogic.scala 711:122]
  wire [2:0] _GEN_1273 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 ?
    _GEN_1263 : _GEN_1269; // @[\\src\\main\\scala\\GameLogic.scala 711:122]
  wire  _GEN_1274 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 | _GEN_1266; // @[\\src\\main\\scala\\GameLogic.scala 711:122 699:31]
  wire  _GEN_1275 = $signed(spriteXRegs_3) > 11'sh113 & $signed(spriteXRegs_3) < 11'sh133 & _T_815 & _T_817 ? 1'h0 :
    _T_832; // @[\\src\\main\\scala\\GameLogic.scala 711:122 700:31]
  wire  _GEN_1276 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 702:116 695:30 703:32]
  wire [1:0] _GEN_1278 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3)
     > 10'sh12c & $signed(spriteYRegs_3) < 10'sh14c ? _GEN_1262 : _GEN_1272; // @[\\src\\main\\scala\\GameLogic.scala 702:116]
  wire [2:0] _GEN_1279 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3)
     > 10'sh12c & $signed(spriteYRegs_3) < 10'sh14c ? _GEN_1263 : _GEN_1273; // @[\\src\\main\\scala\\GameLogic.scala 702:116]
  wire  _GEN_1280 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c | _GEN_1270; // @[\\src\\main\\scala\\GameLogic.scala 702:116 697:30]
  wire  _GEN_1281 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c ? 1'h0 : _T_825; // @[\\src\\main\\scala\\GameLogic.scala 702:116 698:31]
  wire  _GEN_1282 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c | _GEN_1274; // @[\\src\\main\\scala\\GameLogic.scala 702:116 699:31]
  wire  _GEN_1283 = $signed(spriteXRegs_3) > 11'she3 & $signed(spriteXRegs_3) < 11'sh103 & $signed(spriteYRegs_3) > 10'sh12c
     & $signed(spriteYRegs_3) < 10'sh14c ? 1'h0 : _GEN_1275; // @[\\src\\main\\scala\\GameLogic.scala 702:116 700:31]
  wire [2:0] _GEN_1284 = _T ? 3'h4 : _GEN_1279; // @[\\src\\main\\scala\\GameLogic.scala 690:28 691:18]
  wire  _GEN_1285 = _T ? spriteVisibleRegs_3 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 690:28 125:34 694:30]
  wire  _GEN_1286 = _T ? spriteVisibleRegs_7 : _GEN_1276; // @[\\src\\main\\scala\\GameLogic.scala 690:28 125:34]
  wire  _GEN_1287 = _T ? spriteVisibleRegs_8 : _T_818; // @[\\src\\main\\scala\\GameLogic.scala 690:28 125:34]
  wire  _GEN_1288 = _T ? spriteVisibleRegs_9 : _GEN_1280; // @[\\src\\main\\scala\\GameLogic.scala 690:28 125:34]
  wire  _GEN_1289 = _T ? spriteVisibleRegs_10 : _GEN_1281; // @[\\src\\main\\scala\\GameLogic.scala 690:28 125:34]
  wire  _GEN_1290 = _T ? spriteVisibleRegs_11 : _GEN_1282; // @[\\src\\main\\scala\\GameLogic.scala 690:28 125:34]
  wire  _GEN_1291 = _T ? spriteVisibleRegs_12 : _GEN_1283; // @[\\src\\main\\scala\\GameLogic.scala 690:28 125:34]
  wire [1:0] _GEN_1292 = _T ? lvlReg : _GEN_1278; // @[\\src\\main\\scala\\GameLogic.scala 211:23 690:28]
  wire [9:0] _GEN_1293 = _T_83 ? 10'h280 : viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 758:34 759:21 201:28]
  wire [8:0] _GEN_1294 = _T_83 ? 9'h1e0 : viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 758:34 760:21 202:28]
  wire [9:0] _GEN_1295 = _T_76 ? 10'h0 : _GEN_1293; // @[\\src\\main\\scala\\GameLogic.scala 755:34 756:21]
  wire [8:0] _GEN_1296 = _T_76 ? 9'h1e0 : _GEN_1294; // @[\\src\\main\\scala\\GameLogic.scala 755:34 757:21]
  wire [9:0] _GEN_1297 = _T_69 ? 10'h280 : _GEN_1295; // @[\\src\\main\\scala\\GameLogic.scala 752:28 753:21]
  wire [8:0] _GEN_1298 = _T_69 ? 9'h0 : _GEN_1296; // @[\\src\\main\\scala\\GameLogic.scala 752:28 754:21]
  wire [9:0] _spriteYRegs_14_T_2 = $signed(spriteYRegs_14) + 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 770:48]
  wire [9:0] _GEN_1299 = $signed(spriteYRegs_14) < 10'sh1c0 ? $signed(_spriteYRegs_14_T_2) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 769:48 770:29]
  wire [9:0] _spriteYRegs_14_T_5 = $signed(spriteYRegs_14) - 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 774:48]
  wire [9:0] _GEN_1300 = $signed(spriteYRegs_14) > 10'sh20 ? $signed(_spriteYRegs_14_T_5) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 773:40 774:29]
  wire [9:0] _GEN_1301 = io_btnU ? $signed(_GEN_1300) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 772:29]
  wire [9:0] _GEN_1302 = io_btnD ? $signed(_GEN_1299) : $signed(_GEN_1301); // @[\\src\\main\\scala\\GameLogic.scala 768:23]
  wire [9:0] _spriteYRegs_3_T_2 = $signed(spriteYRegs_3) + 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 314:58]
  wire [9:0] _GEN_1303 = $signed(spriteYRegs_3) < 10'sh1c0 ? $signed(_spriteYRegs_3_T_2) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 313:51 314:32]
  wire [9:0] _spriteYRegs_3_T_5 = $signed(spriteYRegs_3) - 10'sh2; // @[\\src\\main\\scala\\GameLogic.scala 318:58]
  wire [9:0] _GEN_1304 = $signed(spriteYRegs_3) > 10'sh20 ? $signed(_spriteYRegs_3_T_5) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 317:43 318:32]
  wire [9:0] _GEN_1305 = io_btnU ? $signed(_GEN_1304) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 316:25]
  wire [9:0] _GEN_1306 = io_btnD ? $signed(_GEN_1303) : $signed(_GEN_1305); // @[\\src\\main\\scala\\GameLogic.scala 312:19]
  wire [10:0] _spriteXRegs_3_T_2 = $signed(spriteXRegs_3) + 11'sh2; // @[\\src\\main\\scala\\GameLogic.scala 323:58]
  wire [10:0] _GEN_1307 = $signed(spriteXRegs_3) < 11'sh260 ? $signed(_spriteXRegs_3_T_2) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 322:51 323:32]
  wire [10:0] _spriteXRegs_3_T_5 = $signed(spriteXRegs_3) - 11'sh2; // @[\\src\\main\\scala\\GameLogic.scala 327:58]
  wire [10:0] _GEN_1308 = $signed(spriteXRegs_3) > 11'sh20 ? $signed(_spriteXRegs_3_T_5) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 326:43 327:32]
  wire [10:0] _GEN_1309 = io_btnL ? $signed(_GEN_1308) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 325:25]
  wire [10:0] _GEN_1310 = io_btnR ? $signed(_GEN_1307) : $signed(_GEN_1309); // @[\\src\\main\\scala\\GameLogic.scala 321:19]
  wire [9:0] _GEN_1311 = _T ? $signed(_GEN_1302) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 767:28]
  wire [9:0] _GEN_1312 = _T ? $signed(_GEN_1) : $signed(_GEN_1306); // @[\\src\\main\\scala\\GameLogic.scala 767:28]
  wire [10:0] _GEN_1313 = _T ? $signed(_GEN_0) : $signed(_GEN_1310); // @[\\src\\main\\scala\\GameLogic.scala 767:28]
  wire [2:0] _GEN_1314 = _T_5 ? 3'h6 : 3'h5; // @[\\src\\main\\scala\\GameLogic.scala 782:30 783:18 785:18]
  wire  _cursorOnReturn_T_3 = $signed(spriteYRegs_3) >= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 801:24]
  wire  _cursorOnReturn_T_4 = $signed(spriteXRegs_3) >= 11'sh110 & $signed(spriteXRegs_3) <= 11'sh170 &
    _cursorOnReturn_T_3; // @[\\src\\main\\scala\\GameLogic.scala 800:79]
  wire  cursorOnReturn = _cursorOnReturn_T_4 & $signed(spriteYRegs_3) <= 10'sh124; // @[\\src\\main\\scala\\GameLogic.scala 801:33]
  wire  _spriteVisibleRegs_52_T = ~cursorOnReturn; // @[\\src\\main\\scala\\GameLogic.scala 803:32]
  wire  _GEN_1323 = cursorOnReturn & io_btnC | gameOverReturnPressed; // @[\\src\\main\\scala\\GameLogic.scala 815:39 816:31 247:38]
  wire [2:0] _GEN_1325 = 3'h5 == stateReg ? 3'h0 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 336:20 823:16 113:25]
  wire  _GEN_1326 = 3'h6 == stateReg ? 1'h0 : spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 336:20 790:29 125:34]
  wire  _GEN_1327 = 3'h6 == stateReg | spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 336:20 793:29 125:34]
  wire  _GEN_1328 = 3'h6 == stateReg | spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 336:20 794:29 125:34]
  wire  _GEN_1329 = 3'h6 == stateReg | spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 336:20 795:29 125:34]
  wire  _GEN_1330 = 3'h6 == stateReg | spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 336:20 796:29 125:34]
  wire  _GEN_1331 = 3'h6 == stateReg | spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 336:20 797:29 125:34]
  wire  _GEN_1332 = 3'h6 == stateReg | spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 336:20 798:29 125:34]
  wire  _GEN_1333 = 3'h6 == stateReg ? ~cursorOnReturn : spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 336:20 803:29 125:34]
  wire  _GEN_1334 = 3'h6 == stateReg ? _spriteVisibleRegs_52_T : spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 336:20 804:29 125:34]
  wire  _GEN_1335 = 3'h6 == stateReg ? _spriteVisibleRegs_52_T : spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 336:20 805:29 125:34]
  wire  _GEN_1336 = 3'h6 == stateReg ? cursorOnReturn : spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 336:20 806:29 125:34]
  wire  _GEN_1337 = 3'h6 == stateReg ? cursorOnReturn : spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 336:20 807:29 125:34]
  wire  _GEN_1338 = 3'h6 == stateReg ? cursorOnReturn : spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 336:20 808:29 125:34]
  wire  _GEN_1339 = 3'h6 == stateReg | spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 336:20 811:28 125:34]
  wire [9:0] _GEN_1340 = 3'h6 == stateReg ? $signed(_GEN_1306) : $signed(_GEN_1); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [10:0] _GEN_1341 = 3'h6 == stateReg ? $signed(_GEN_1310) : $signed(_GEN_0); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1342 = 3'h6 == stateReg ? _GEN_1323 : gameOverReturnPressed; // @[\\src\\main\\scala\\GameLogic.scala 336:20 247:38]
  wire [2:0] _GEN_1343 = 3'h6 == stateReg ? 3'h5 : _GEN_1325; // @[\\src\\main\\scala\\GameLogic.scala 336:20 819:16]
  wire  _GEN_1344 = 3'h6 == stateReg ? 1'h0 : 3'h5 == stateReg; // @[\\src\\main\\scala\\GameLogic.scala 336:20 100:22]
  wire [9:0] _GEN_1345 = 3'h4 == stateReg ? $signed(_GEN_1311) : $signed(_GEN_17); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [9:0] _GEN_1346 = 3'h4 == stateReg ? $signed(_GEN_1312) : $signed(_GEN_1340); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [10:0] _GEN_1347 = 3'h4 == stateReg ? $signed(_GEN_1313) : $signed(_GEN_1341); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [2:0] _GEN_1348 = 3'h4 == stateReg ? _GEN_1314 : _GEN_1343; // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1349 = 3'h4 == stateReg ? spriteVisibleRegs_14 : _GEN_1326; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1350 = 3'h4 == stateReg ? spriteVisibleRegs_46 : _GEN_1327; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1351 = 3'h4 == stateReg ? spriteVisibleRegs_47 : _GEN_1328; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1352 = 3'h4 == stateReg ? spriteVisibleRegs_48 : _GEN_1329; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1353 = 3'h4 == stateReg ? spriteVisibleRegs_49 : _GEN_1330; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1354 = 3'h4 == stateReg ? spriteVisibleRegs_50 : _GEN_1331; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1355 = 3'h4 == stateReg ? spriteVisibleRegs_51 : _GEN_1332; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1356 = 3'h4 == stateReg ? spriteVisibleRegs_52 : _GEN_1333; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1357 = 3'h4 == stateReg ? spriteVisibleRegs_53 : _GEN_1334; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1358 = 3'h4 == stateReg ? spriteVisibleRegs_54 : _GEN_1335; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1359 = 3'h4 == stateReg ? spriteVisibleRegs_55 : _GEN_1336; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1360 = 3'h4 == stateReg ? spriteVisibleRegs_56 : _GEN_1337; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1361 = 3'h4 == stateReg ? spriteVisibleRegs_57 : _GEN_1338; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1362 = 3'h4 == stateReg ? spriteVisibleRegs_3 : _GEN_1339; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1363 = 3'h4 == stateReg ? gameOverReturnPressed : _GEN_1342; // @[\\src\\main\\scala\\GameLogic.scala 336:20 247:38]
  wire  _GEN_1364 = 3'h4 == stateReg ? 1'h0 : _GEN_1344; // @[\\src\\main\\scala\\GameLogic.scala 336:20 100:22]
  wire [5:0] _GEN_1365 = 3'h3 == stateReg ? 6'h0 : nextSpriteToSpawn; // @[\\src\\main\\scala\\GameLogic.scala 336:20 736:25 232:34]
  wire [7:0] _GEN_1366 = 3'h3 == stateReg ? 8'h0 : spawnDelayCounter; // @[\\src\\main\\scala\\GameLogic.scala 336:20 737:25 231:34]
  wire [10:0] _GEN_1367 = 3'h3 == stateReg ? $signed(11'sh260) : $signed(_GEN_16); // @[\\src\\main\\scala\\GameLogic.scala 336:20 739:23]
  wire [9:0] _GEN_1368 = 3'h3 == stateReg ? $signed(10'sh140) : $signed(_GEN_1345); // @[\\src\\main\\scala\\GameLogic.scala 336:20 740:23]
  wire  _GEN_1369 = 3'h3 == stateReg ? 1'h0 : _GEN_1362; // @[\\src\\main\\scala\\GameLogic.scala 336:20 741:28]
  wire  _GEN_1370 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 336:20 742:28 125:34]
  wire  _GEN_1371 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 336:20 743:28 125:34]
  wire  _GEN_1372 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 336:20 744:28 125:34]
  wire  _GEN_1373 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 336:20 745:29 125:34]
  wire  _GEN_1374 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 336:20 746:29 125:34]
  wire  _GEN_1375 = 3'h3 == stateReg ? 1'h0 : spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 336:20 747:29 125:34]
  wire  _GEN_1376 = 3'h3 == stateReg | _GEN_1349; // @[\\src\\main\\scala\\GameLogic.scala 336:20 748:29]
  wire  _GEN_1377 = 3'h3 == stateReg | _GEN_123; // @[\\src\\main\\scala\\GameLogic.scala 336:20 749:29]
  wire  _GEN_1378 = 3'h3 == stateReg | _GEN_124; // @[\\src\\main\\scala\\GameLogic.scala 336:20 750:29]
  wire  _GEN_1379 = 3'h3 == stateReg | _GEN_125; // @[\\src\\main\\scala\\GameLogic.scala 336:20 751:29]
  wire [9:0] _GEN_1380 = 3'h3 == stateReg ? _GEN_1297 : viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 336:20 201:28]
  wire [8:0] _GEN_1381 = 3'h3 == stateReg ? _GEN_1298 : viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 336:20 202:28]
  wire [2:0] _GEN_1382 = 3'h3 == stateReg ? 3'h4 : _GEN_1348; // @[\\src\\main\\scala\\GameLogic.scala 336:20 762:16]
  wire [9:0] _GEN_1383 = 3'h3 == stateReg ? $signed(_GEN_1) : $signed(_GEN_1346); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [10:0] _GEN_1384 = 3'h3 == stateReg ? $signed(_GEN_0) : $signed(_GEN_1347); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1385 = 3'h3 == stateReg ? spriteVisibleRegs_46 : _GEN_1350; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1386 = 3'h3 == stateReg ? spriteVisibleRegs_47 : _GEN_1351; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1387 = 3'h3 == stateReg ? spriteVisibleRegs_48 : _GEN_1352; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1388 = 3'h3 == stateReg ? spriteVisibleRegs_49 : _GEN_1353; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1389 = 3'h3 == stateReg ? spriteVisibleRegs_50 : _GEN_1354; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1390 = 3'h3 == stateReg ? spriteVisibleRegs_51 : _GEN_1355; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1391 = 3'h3 == stateReg ? spriteVisibleRegs_52 : _GEN_1356; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1392 = 3'h3 == stateReg ? spriteVisibleRegs_53 : _GEN_1357; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1393 = 3'h3 == stateReg ? spriteVisibleRegs_54 : _GEN_1358; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1394 = 3'h3 == stateReg ? spriteVisibleRegs_55 : _GEN_1359; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1395 = 3'h3 == stateReg ? spriteVisibleRegs_56 : _GEN_1360; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1396 = 3'h3 == stateReg ? spriteVisibleRegs_57 : _GEN_1361; // @[\\src\\main\\scala\\GameLogic.scala 336:20 125:34]
  wire  _GEN_1397 = 3'h3 == stateReg ? gameOverReturnPressed : _GEN_1363; // @[\\src\\main\\scala\\GameLogic.scala 336:20 247:38]
  wire  _GEN_1398 = 3'h3 == stateReg ? 1'h0 : _GEN_1364; // @[\\src\\main\\scala\\GameLogic.scala 336:20 100:22]
  wire  _GEN_1433 = 3'h2 == stateReg ? 1'h0 : _GEN_1398; // @[\\src\\main\\scala\\GameLogic.scala 336:20 100:22]
  wire [26:0] _GEN_1436 = 3'h1 == stateReg ? $signed(_GEN_399) : $signed({{16{_GEN_18[10]}},_GEN_18}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1439 = 3'h1 == stateReg ? _GEN_402 : spriteScaleTypeRegs_0; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1441 = 3'h1 == stateReg ? $signed(_GEN_404) : $signed({{16{_GEN_20[10]}},_GEN_20}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1444 = 3'h1 == stateReg ? _GEN_407 : spriteScaleTypeRegs_1; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1446 = 3'h1 == stateReg ? $signed(_GEN_409) : $signed({{16{_GEN_22[10]}},_GEN_22}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1449 = 3'h1 == stateReg ? _GEN_412 : spriteScaleTypeRegs_2; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1451 = 3'h1 == stateReg ? $signed(_GEN_414) : $signed({{16{_GEN_24[10]}},_GEN_24}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1454 = 3'h1 == stateReg ? _GEN_417 : spriteScaleTypeRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1456 = 3'h1 == stateReg ? $signed(_GEN_419) : $signed({{16{_GEN_26[10]}},_GEN_26}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1459 = 3'h1 == stateReg ? _GEN_422 : spriteScaleTypeRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1461 = 3'h1 == stateReg ? $signed(_GEN_424) : $signed({{16{_GEN_28[10]}},_GEN_28}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1464 = 3'h1 == stateReg ? _GEN_427 : spriteScaleTypeRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1466 = 3'h1 == stateReg ? $signed(_GEN_429) : $signed({{16{_GEN_30[10]}},_GEN_30}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1469 = 3'h1 == stateReg ? _GEN_432 : spriteScaleTypeRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1471 = 3'h1 == stateReg ? $signed(_GEN_434) : $signed({{16{_GEN_32[10]}},_GEN_32}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1474 = 3'h1 == stateReg ? _GEN_437 : spriteScaleTypeRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1476 = 3'h1 == stateReg ? $signed(_GEN_439) : $signed({{16{_GEN_34[10]}},_GEN_34}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1479 = 3'h1 == stateReg ? _GEN_442 : spriteScaleTypeRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1481 = 3'h1 == stateReg ? $signed(_GEN_444) : $signed({{16{_GEN_36[10]}},_GEN_36}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1484 = 3'h1 == stateReg ? _GEN_447 : spriteScaleTypeRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  wire [26:0] _GEN_1486 = 3'h1 == stateReg ? $signed(_GEN_449) : $signed({{16{_GEN_38[10]}},_GEN_38}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1490 = 3'h1 == stateReg ? $signed(_GEN_453) : $signed({{16{_GEN_40[10]}},_GEN_40}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1494 = 3'h1 == stateReg ? $signed(_GEN_457) : $signed({{16{_GEN_42[10]}},_GEN_42}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1498 = 3'h1 == stateReg ? $signed(_GEN_461) : $signed({{16{_GEN_44[10]}},_GEN_44}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1502 = 3'h1 == stateReg ? $signed(_GEN_465) : $signed({{16{_GEN_46[10]}},_GEN_46}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1506 = 3'h1 == stateReg ? $signed(_GEN_469) : $signed({{16{_GEN_48[10]}},_GEN_48}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1510 = 3'h1 == stateReg ? $signed(_GEN_473) : $signed({{16{_GEN_50[10]}},_GEN_50}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1514 = 3'h1 == stateReg ? $signed(_GEN_477) : $signed({{16{_GEN_52[10]}},_GEN_52}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1518 = 3'h1 == stateReg ? $signed(_GEN_481) : $signed({{16{_GEN_54[10]}},_GEN_54}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1522 = 3'h1 == stateReg ? $signed(_GEN_485) : $signed({{16{_GEN_56[10]}},_GEN_56}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1526 = 3'h1 == stateReg ? $signed(_GEN_489) : $signed({{16{_GEN_58[10]}},_GEN_58}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1530 = 3'h1 == stateReg ? $signed(_GEN_493) : $signed({{16{_GEN_60[10]}},_GEN_60}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1534 = 3'h1 == stateReg ? $signed(_GEN_497) : $signed({{16{_GEN_62[10]}},_GEN_62}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1538 = 3'h1 == stateReg ? $signed(_GEN_501) : $signed({{16{_GEN_64[10]}},_GEN_64}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1542 = 3'h1 == stateReg ? $signed(_GEN_505) : $signed({{16{_GEN_66[10]}},_GEN_66}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1546 = 3'h1 == stateReg ? $signed(_GEN_509) : $signed({{16{_GEN_68[10]}},_GEN_68}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1550 = 3'h1 == stateReg ? $signed(_GEN_513) : $signed({{16{_GEN_70[10]}},_GEN_70}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1554 = 3'h1 == stateReg ? $signed(_GEN_517) : $signed({{16{_GEN_72[10]}},_GEN_72}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1558 = 3'h1 == stateReg ? $signed(_GEN_521) : $signed({{16{_GEN_74[10]}},_GEN_74}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1562 = 3'h1 == stateReg ? $signed(_GEN_525) : $signed({{16{_GEN_76[10]}},_GEN_76}); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire  _GEN_1662 = 3'h1 == stateReg ? 1'h0 : _GEN_1433; // @[\\src\\main\\scala\\GameLogic.scala 336:20 100:22]
  wire  _GEN_1674 = 3'h0 == stateReg ? _GEN_196 : _GEN_114; // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1722 = 3'h0 == stateReg ? $signed({{16{_GEN_18[10]}},_GEN_18}) : $signed(_GEN_1436); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1727 = 3'h0 == stateReg ? $signed({{16{_GEN_20[10]}},_GEN_20}) : $signed(_GEN_1441); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1732 = 3'h0 == stateReg ? $signed({{16{_GEN_22[10]}},_GEN_22}) : $signed(_GEN_1446); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1737 = 3'h0 == stateReg ? $signed({{16{_GEN_24[10]}},_GEN_24}) : $signed(_GEN_1451); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1742 = 3'h0 == stateReg ? $signed({{16{_GEN_26[10]}},_GEN_26}) : $signed(_GEN_1456); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1747 = 3'h0 == stateReg ? $signed({{16{_GEN_28[10]}},_GEN_28}) : $signed(_GEN_1461); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1752 = 3'h0 == stateReg ? $signed({{16{_GEN_30[10]}},_GEN_30}) : $signed(_GEN_1466); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1757 = 3'h0 == stateReg ? $signed({{16{_GEN_32[10]}},_GEN_32}) : $signed(_GEN_1471); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1762 = 3'h0 == stateReg ? $signed({{16{_GEN_34[10]}},_GEN_34}) : $signed(_GEN_1476); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1767 = 3'h0 == stateReg ? $signed({{16{_GEN_36[10]}},_GEN_36}) : $signed(_GEN_1481); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1772 = 3'h0 == stateReg ? $signed({{16{_GEN_38[10]}},_GEN_38}) : $signed(_GEN_1486); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1776 = 3'h0 == stateReg ? $signed({{16{_GEN_40[10]}},_GEN_40}) : $signed(_GEN_1490); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1780 = 3'h0 == stateReg ? $signed({{16{_GEN_42[10]}},_GEN_42}) : $signed(_GEN_1494); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1784 = 3'h0 == stateReg ? $signed({{16{_GEN_44[10]}},_GEN_44}) : $signed(_GEN_1498); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1788 = 3'h0 == stateReg ? $signed({{16{_GEN_46[10]}},_GEN_46}) : $signed(_GEN_1502); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1792 = 3'h0 == stateReg ? $signed({{16{_GEN_48[10]}},_GEN_48}) : $signed(_GEN_1506); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1796 = 3'h0 == stateReg ? $signed({{16{_GEN_50[10]}},_GEN_50}) : $signed(_GEN_1510); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1800 = 3'h0 == stateReg ? $signed({{16{_GEN_52[10]}},_GEN_52}) : $signed(_GEN_1514); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1804 = 3'h0 == stateReg ? $signed({{16{_GEN_54[10]}},_GEN_54}) : $signed(_GEN_1518); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1808 = 3'h0 == stateReg ? $signed({{16{_GEN_56[10]}},_GEN_56}) : $signed(_GEN_1522); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1812 = 3'h0 == stateReg ? $signed({{16{_GEN_58[10]}},_GEN_58}) : $signed(_GEN_1526); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1816 = 3'h0 == stateReg ? $signed({{16{_GEN_60[10]}},_GEN_60}) : $signed(_GEN_1530); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1820 = 3'h0 == stateReg ? $signed({{16{_GEN_62[10]}},_GEN_62}) : $signed(_GEN_1534); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1824 = 3'h0 == stateReg ? $signed({{16{_GEN_64[10]}},_GEN_64}) : $signed(_GEN_1538); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1828 = 3'h0 == stateReg ? $signed({{16{_GEN_66[10]}},_GEN_66}) : $signed(_GEN_1542); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1832 = 3'h0 == stateReg ? $signed({{16{_GEN_68[10]}},_GEN_68}) : $signed(_GEN_1546); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1836 = 3'h0 == stateReg ? $signed({{16{_GEN_70[10]}},_GEN_70}) : $signed(_GEN_1550); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1840 = 3'h0 == stateReg ? $signed({{16{_GEN_72[10]}},_GEN_72}) : $signed(_GEN_1554); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1844 = 3'h0 == stateReg ? $signed({{16{_GEN_74[10]}},_GEN_74}) : $signed(_GEN_1558); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_1848 = 3'h0 == stateReg ? $signed({{16{_GEN_76[10]}},_GEN_76}) : $signed(_GEN_1562); // @[\\src\\main\\scala\\GameLogic.scala 336:20]
  wire [26:0] _GEN_2091 = reset ? $signed(27'sh0) : $signed(_GEN_1722); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2093 = reset ? $signed(27'sh0) : $signed(_GEN_1727); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2095 = reset ? $signed(27'sh0) : $signed(_GEN_1732); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2097 = reset ? $signed(27'sh0) : $signed(_GEN_1737); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2099 = reset ? $signed(27'sh0) : $signed(_GEN_1742); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2101 = reset ? $signed(27'sh0) : $signed(_GEN_1747); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2103 = reset ? $signed(27'sh0) : $signed(_GEN_1752); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2105 = reset ? $signed(27'sh0) : $signed(_GEN_1757); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2107 = reset ? $signed(27'sh0) : $signed(_GEN_1762); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2109 = reset ? $signed(27'sh0) : $signed(_GEN_1767); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2111 = reset ? $signed(27'sh0) : $signed(_GEN_1772); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2113 = reset ? $signed(27'sh0) : $signed(_GEN_1776); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2115 = reset ? $signed(27'sh0) : $signed(_GEN_1780); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2117 = reset ? $signed(27'sh0) : $signed(_GEN_1784); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2119 = reset ? $signed(27'sh0) : $signed(_GEN_1788); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2121 = reset ? $signed(27'sh0) : $signed(_GEN_1792); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2123 = reset ? $signed(27'sh0) : $signed(_GEN_1796); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2125 = reset ? $signed(27'sh0) : $signed(_GEN_1800); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2127 = reset ? $signed(27'sh0) : $signed(_GEN_1804); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2129 = reset ? $signed(27'sh0) : $signed(_GEN_1808); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2131 = reset ? $signed(27'sh0) : $signed(_GEN_1812); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2133 = reset ? $signed(27'sh0) : $signed(_GEN_1816); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2135 = reset ? $signed(27'sh0) : $signed(_GEN_1820); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2137 = reset ? $signed(27'sh0) : $signed(_GEN_1824); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2139 = reset ? $signed(27'sh0) : $signed(_GEN_1828); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2141 = reset ? $signed(27'sh0) : $signed(_GEN_1832); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2143 = reset ? $signed(27'sh0) : $signed(_GEN_1836); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2145 = reset ? $signed(27'sh0) : $signed(_GEN_1840); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2147 = reset ? $signed(27'sh0) : $signed(_GEN_1844); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  wire [26:0] _GEN_2149 = reset ? $signed(27'sh0) : $signed(_GEN_1848); // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
  Difficulty difficulty ( // @[\\src\\main\\scala\\GameLogic.scala 209:26]
    .clock(difficulty_clock),
    .reset(difficulty_reset),
    .io_level(difficulty_io_level),
    .io_speed(difficulty_io_speed),
    .io_resetSpeed(difficulty_io_resetSpeed)
  );
  LFSR lfsr ( // @[\\src\\main\\scala\\GameLogic.scala 250:20]
    .clock(lfsr_clock),
    .reset(lfsr_reset),
    .io_out_0(lfsr_io_out_0),
    .io_out_1(lfsr_io_out_1),
    .io_out_2(lfsr_io_out_2),
    .io_out_3(lfsr_io_out_3),
    .io_out_4(lfsr_io_out_4),
    .io_out_5(lfsr_io_out_5),
    .io_out_6(lfsr_io_out_6),
    .io_out_7(lfsr_io_out_7),
    .io_out_8(lfsr_io_out_8),
    .io_out_9(lfsr_io_out_9),
    .io_out_10(lfsr_io_out_10),
    .io_out_11(lfsr_io_out_11),
    .io_out_12(lfsr_io_out_12),
    .io_out_13(lfsr_io_out_13),
    .io_out_14(lfsr_io_out_14),
    .io_out_15(lfsr_io_out_15),
    .io_out_16(lfsr_io_out_16),
    .io_out_17(lfsr_io_out_17),
    .io_out_18(lfsr_io_out_18),
    .io_out_19(lfsr_io_out_19),
    .io_out_20(lfsr_io_out_20),
    .io_out_21(lfsr_io_out_21),
    .io_out_22(lfsr_io_out_22),
    .io_out_23(lfsr_io_out_23),
    .io_out_24(lfsr_io_out_24),
    .io_out_25(lfsr_io_out_25),
    .io_out_26(lfsr_io_out_26),
    .io_out_27(lfsr_io_out_27),
    .io_out_28(lfsr_io_out_28),
    .io_out_29(lfsr_io_out_29)
  );
  assign io_spriteXPosition_3 = spriteXRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_7 = spriteXRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_8 = spriteXRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_9 = spriteXRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_10 = spriteXRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_11 = spriteXRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_12 = spriteXRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_13 = spriteXRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_14 = spriteXRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_16 = spriteXRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_17 = spriteXRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_18 = spriteXRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_19 = spriteXRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_20 = spriteXRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_21 = spriteXRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_22 = spriteXRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_23 = spriteXRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_24 = spriteXRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_25 = spriteXRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_26 = spriteXRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_27 = spriteXRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_28 = spriteXRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_29 = spriteXRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_30 = spriteXRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_31 = spriteXRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_32 = spriteXRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_33 = spriteXRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_34 = spriteXRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_35 = spriteXRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_36 = spriteXRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_37 = spriteXRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_38 = spriteXRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_39 = spriteXRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_40 = spriteXRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_41 = spriteXRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_42 = spriteXRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_43 = spriteXRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_44 = spriteXRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_45 = spriteXRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_46 = spriteXRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_47 = spriteXRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_48 = spriteXRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_49 = spriteXRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_50 = spriteXRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_51 = spriteXRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_52 = spriteXRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_53 = spriteXRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_54 = spriteXRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_55 = spriteXRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_56 = spriteXRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_57 = spriteXRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_58 = spriteXRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_59 = spriteXRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_60 = spriteXRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_61 = spriteXRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_62 = spriteXRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteXPosition_63 = spriteXRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 180:27]
  assign io_spriteYPosition_3 = spriteYRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_7 = spriteYRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_8 = spriteYRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_9 = spriteYRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_10 = spriteYRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_11 = spriteYRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_12 = spriteYRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_13 = spriteYRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_14 = spriteYRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_16 = spriteYRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_17 = spriteYRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_18 = spriteYRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_19 = spriteYRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_20 = spriteYRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_21 = spriteYRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_22 = spriteYRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_23 = spriteYRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_24 = spriteYRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_25 = spriteYRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_26 = spriteYRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_27 = spriteYRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_28 = spriteYRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_29 = spriteYRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_30 = spriteYRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_31 = spriteYRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_32 = spriteYRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_33 = spriteYRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_34 = spriteYRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_35 = spriteYRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_36 = spriteYRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_37 = spriteYRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_38 = spriteYRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_39 = spriteYRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_40 = spriteYRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_41 = spriteYRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_42 = spriteYRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_43 = spriteYRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_44 = spriteYRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_45 = spriteYRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_46 = spriteYRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_47 = spriteYRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_48 = spriteYRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_49 = spriteYRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_50 = spriteYRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_51 = spriteYRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_52 = spriteYRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_53 = spriteYRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_54 = spriteYRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_55 = spriteYRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_56 = spriteYRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_57 = spriteYRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_58 = spriteYRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_59 = spriteYRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_60 = spriteYRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_61 = spriteYRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_62 = spriteYRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteYPosition_63 = spriteYRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 181:27]
  assign io_spriteVisible_3 = spriteVisibleRegs_3; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_4 = spriteVisibleRegs_4; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_5 = spriteVisibleRegs_5; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_6 = spriteVisibleRegs_6; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_7 = spriteVisibleRegs_7; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_8 = spriteVisibleRegs_8; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_9 = spriteVisibleRegs_9; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_10 = spriteVisibleRegs_10; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_11 = spriteVisibleRegs_11; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_12 = spriteVisibleRegs_12; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_13 = spriteVisibleRegs_13; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_14 = spriteVisibleRegs_14; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_15 = spriteVisibleRegs_15; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_16 = spriteVisibleRegs_16; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_17 = spriteVisibleRegs_17; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_18 = spriteVisibleRegs_18; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_19 = spriteVisibleRegs_19; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_20 = spriteVisibleRegs_20; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_21 = spriteVisibleRegs_21; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_22 = spriteVisibleRegs_22; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_23 = spriteVisibleRegs_23; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_24 = spriteVisibleRegs_24; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_25 = spriteVisibleRegs_25; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_26 = spriteVisibleRegs_26; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_27 = spriteVisibleRegs_27; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_28 = spriteVisibleRegs_28; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_29 = spriteVisibleRegs_29; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_30 = spriteVisibleRegs_30; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_31 = spriteVisibleRegs_31; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_32 = spriteVisibleRegs_32; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_33 = spriteVisibleRegs_33; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_34 = spriteVisibleRegs_34; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_35 = spriteVisibleRegs_35; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_36 = spriteVisibleRegs_36; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_37 = spriteVisibleRegs_37; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_38 = spriteVisibleRegs_38; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_39 = spriteVisibleRegs_39; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_40 = spriteVisibleRegs_40; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_41 = spriteVisibleRegs_41; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_42 = spriteVisibleRegs_42; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_43 = spriteVisibleRegs_43; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_44 = spriteVisibleRegs_44; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_45 = spriteVisibleRegs_45; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_46 = spriteVisibleRegs_46; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_47 = spriteVisibleRegs_47; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_48 = spriteVisibleRegs_48; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_49 = spriteVisibleRegs_49; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_50 = spriteVisibleRegs_50; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_51 = spriteVisibleRegs_51; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_52 = spriteVisibleRegs_52; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_53 = spriteVisibleRegs_53; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_54 = spriteVisibleRegs_54; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_55 = spriteVisibleRegs_55; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_56 = spriteVisibleRegs_56; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_57 = spriteVisibleRegs_57; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_58 = spriteVisibleRegs_58; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_59 = spriteVisibleRegs_59; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_60 = spriteVisibleRegs_60; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_61 = spriteVisibleRegs_61; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_62 = spriteVisibleRegs_62; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteVisible_63 = spriteVisibleRegs_63; // @[\\src\\main\\scala\\GameLogic.scala 177:25]
  assign io_spriteScaleUpHorizontal_16 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1439; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_17 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1444; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_18 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1449; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_19 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1454; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_20 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1459; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_21 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1464; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_22 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1469; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_23 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1474; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_24 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1479; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_25 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1484; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_26 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1439; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_27 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1444; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_28 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1449; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_29 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1454; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_30 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1459; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_31 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1464; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_32 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1469; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_33 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1474; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_34 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1479; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_35 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1484; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_36 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1439; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_37 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1444; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_38 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1449; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_39 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1454; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_40 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1459; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_41 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1464; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_42 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1469; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_43 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1474; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_44 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1479; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_45 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1484; // @[\\src\\main\\scala\\GameLogic.scala 336:20 187:35]
  assign io_spriteScaleUpHorizontal_58 = sprite58ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 193:34]
  assign io_spriteScaleUpHorizontal_59 = sprite59ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 195:34]
  assign io_spriteScaleUpHorizontal_60 = sprite60ScaleUpHorizontal; // @[\\src\\main\\scala\\GameLogic.scala 197:34]
  assign io_spriteScaleUpVertical_16 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1439; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_17 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1444; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_18 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1449; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_19 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1454; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_20 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1459; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_21 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1464; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_22 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1469; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_23 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1474; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_24 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1479; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_25 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1484; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_26 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1439; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_27 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1444; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_28 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1449; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_29 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1454; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_30 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1459; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_31 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1464; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_32 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1469; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_33 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1474; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_34 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1479; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_35 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1484; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_36 = 3'h0 == stateReg ? spriteScaleTypeRegs_0 : _GEN_1439; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_37 = 3'h0 == stateReg ? spriteScaleTypeRegs_1 : _GEN_1444; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_38 = 3'h0 == stateReg ? spriteScaleTypeRegs_2 : _GEN_1449; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_39 = 3'h0 == stateReg ? spriteScaleTypeRegs_3 : _GEN_1454; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_40 = 3'h0 == stateReg ? spriteScaleTypeRegs_4 : _GEN_1459; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_41 = 3'h0 == stateReg ? spriteScaleTypeRegs_5 : _GEN_1464; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_42 = 3'h0 == stateReg ? spriteScaleTypeRegs_6 : _GEN_1469; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_43 = 3'h0 == stateReg ? spriteScaleTypeRegs_7 : _GEN_1474; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_44 = 3'h0 == stateReg ? spriteScaleTypeRegs_8 : _GEN_1479; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_45 = 3'h0 == stateReg ? spriteScaleTypeRegs_9 : _GEN_1484; // @[\\src\\main\\scala\\GameLogic.scala 336:20 188:33]
  assign io_spriteScaleUpVertical_58 = sprite58ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 194:32]
  assign io_spriteScaleUpVertical_59 = sprite59ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 196:32]
  assign io_spriteScaleUpVertical_60 = sprite60ScaleUpVertical; // @[\\src\\main\\scala\\GameLogic.scala 198:32]
  assign io_viewBoxX = viewBoxXReg; // @[\\src\\main\\scala\\GameLogic.scala 205:15]
  assign io_viewBoxY = viewBoxYReg; // @[\\src\\main\\scala\\GameLogic.scala 206:15]
  assign io_frameUpdateDone = 3'h0 == stateReg ? 1'h0 : _GEN_1662; // @[\\src\\main\\scala\\GameLogic.scala 336:20 100:22]
  assign difficulty_clock = clock;
  assign difficulty_reset = reset;
  assign difficulty_io_level = lvlReg; // @[\\src\\main\\scala\\GameLogic.scala 212:23]
  assign difficulty_io_resetSpeed = stateReg == 3'h2 & livesReg == 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 228:50]
  assign lfsr_clock = clock;
  assign lfsr_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 113:25]
      stateReg <= 3'h0; // @[\\src\\main\\scala\\GameLogic.scala 113:25]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          stateReg <= 3'h2; // @[\\src\\main\\scala\\GameLogic.scala 342:20]
        end else begin
          stateReg <= _GEN_126;
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (livesReg > 3'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 684:28]
        stateReg <= 3'h2; // @[\\src\\main\\scala\\GameLogic.scala 685:18]
      end else begin
        stateReg <= _GEN_1179;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      stateReg <= _GEN_1284;
    end else begin
      stateReg <= _GEN_1382;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_3 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_3 <= _GEN_0;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_3 <= _GEN_0;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_3 <= _GEN_0;
    end else begin
      spriteXRegs_3 <= _GEN_1384;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_7 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_7 <= 11'sh100; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_8 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_8 <= 11'sh100; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_9 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_9 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_10 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_10 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_11 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_11 <= 11'sh160; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_12 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_12 <= 11'sh160; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_13 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_13 <= _GEN_14;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteXRegs_13 <= _GEN_397;
      end else begin
        spriteXRegs_13 <= _GEN_14;
      end
    end else begin
      spriteXRegs_13 <= _GEN_14;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_14 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_14 <= _GEN_16;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_14 <= _GEN_16;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_14 <= _GEN_16;
    end else begin
      spriteXRegs_14 <= _GEN_1367;
    end
    spriteXRegs_16 <= _GEN_2091[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_17 <= _GEN_2093[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_18 <= _GEN_2095[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_19 <= _GEN_2097[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_20 <= _GEN_2099[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_21 <= _GEN_2101[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_22 <= _GEN_2103[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_23 <= _GEN_2105[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_24 <= _GEN_2107[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_25 <= _GEN_2109[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_26 <= _GEN_2111[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_27 <= _GEN_2113[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_28 <= _GEN_2115[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_29 <= _GEN_2117[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_30 <= _GEN_2119[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_31 <= _GEN_2121[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_32 <= _GEN_2123[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_33 <= _GEN_2125[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_34 <= _GEN_2127[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_35 <= _GEN_2129[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_36 <= _GEN_2131[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_37 <= _GEN_2133[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_38 <= _GEN_2135[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_39 <= _GEN_2137[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_40 <= _GEN_2139[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_41 <= _GEN_2141[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_42 <= _GEN_2143[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_43 <= _GEN_2145[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_44 <= _GEN_2147[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    spriteXRegs_45 <= _GEN_2149[10:0]; // @[\\src\\main\\scala\\GameLogic.scala 121:{28,28}]
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_46 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_46 <= 11'she0; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_47 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_47 <= 11'sh100; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_48 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_48 <= 11'sh120; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_49 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_49 <= 11'sh140; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_50 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_50 <= 11'sh160; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_51 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_51 <= 11'sh180; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_52 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_52 <= 11'sh110; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_53 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_53 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_54 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_54 <= 11'sh150; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_55 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_55 <= 11'sh110; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_56 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_56 <= 11'sh130; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_57 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_57 <= 11'sh150; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_58 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_58 <= _GEN_102;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 594:29]
        spriteXRegs_58 <= spriteXRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 595:25]
      end else begin
        spriteXRegs_58 <= _GEN_1241;
      end
    end else begin
      spriteXRegs_58 <= _GEN_102;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_59 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_59 <= _GEN_104;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 594:29]
        spriteXRegs_59 <= spriteXRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 597:25]
      end else begin
        spriteXRegs_59 <= _GEN_1242;
      end
    end else begin
      spriteXRegs_59 <= _GEN_104;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_60 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteXRegs_60 <= _GEN_106;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 594:29]
        spriteXRegs_60 <= spriteXRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 599:25]
      end else begin
        spriteXRegs_60 <= _GEN_1243;
      end
    end else begin
      spriteXRegs_60 <= _GEN_106;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_61 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_61 <= 11'sh14; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_62 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_62 <= 11'sh3c; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 121:28]
      spriteXRegs_63 <= 11'sh0; // @[\\src\\main\\scala\\GameLogic.scala 121:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteXRegs_63 <= 11'sh64; // @[\\src\\main\\scala\\GameLogic.scala 161:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_3 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_3 <= _GEN_1;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_3 <= _GEN_1;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_3 <= _GEN_1;
    end else begin
      spriteYRegs_3 <= _GEN_1383;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_7 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_7 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_8 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_8 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_9 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_9 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_10 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_10 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_11 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_11 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_12 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_12 <= 10'sh12c; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_13 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_13 <= _GEN_15;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_13 <= _GEN_395;
      end else begin
        spriteYRegs_13 <= _GEN_15;
      end
    end else begin
      spriteYRegs_13 <= _GEN_15;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_14 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_14 <= _GEN_17;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_14 <= _GEN_17;
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_14 <= _GEN_17;
    end else begin
      spriteYRegs_14 <= _GEN_1368;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_16 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_16 <= _GEN_19;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_16 <= _GEN_245;
      end else begin
        spriteYRegs_16 <= _GEN_19;
      end
    end else begin
      spriteYRegs_16 <= _GEN_19;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_17 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_17 <= _GEN_21;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_17 <= _GEN_250;
      end else begin
        spriteYRegs_17 <= _GEN_21;
      end
    end else begin
      spriteYRegs_17 <= _GEN_21;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_18 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_18 <= _GEN_23;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_18 <= _GEN_255;
      end else begin
        spriteYRegs_18 <= _GEN_23;
      end
    end else begin
      spriteYRegs_18 <= _GEN_23;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_19 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_19 <= _GEN_25;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_19 <= _GEN_260;
      end else begin
        spriteYRegs_19 <= _GEN_25;
      end
    end else begin
      spriteYRegs_19 <= _GEN_25;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_20 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_20 <= _GEN_27;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_20 <= _GEN_265;
      end else begin
        spriteYRegs_20 <= _GEN_27;
      end
    end else begin
      spriteYRegs_20 <= _GEN_27;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_21 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_21 <= _GEN_29;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_21 <= _GEN_270;
      end else begin
        spriteYRegs_21 <= _GEN_29;
      end
    end else begin
      spriteYRegs_21 <= _GEN_29;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_22 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_22 <= _GEN_31;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_22 <= _GEN_275;
      end else begin
        spriteYRegs_22 <= _GEN_31;
      end
    end else begin
      spriteYRegs_22 <= _GEN_31;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_23 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_23 <= _GEN_33;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_23 <= _GEN_280;
      end else begin
        spriteYRegs_23 <= _GEN_33;
      end
    end else begin
      spriteYRegs_23 <= _GEN_33;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_24 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_24 <= _GEN_35;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_24 <= _GEN_285;
      end else begin
        spriteYRegs_24 <= _GEN_35;
      end
    end else begin
      spriteYRegs_24 <= _GEN_35;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_25 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_25 <= _GEN_37;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_25 <= _GEN_290;
      end else begin
        spriteYRegs_25 <= _GEN_37;
      end
    end else begin
      spriteYRegs_25 <= _GEN_37;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_26 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_26 <= _GEN_39;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_26 <= _GEN_295;
      end else begin
        spriteYRegs_26 <= _GEN_39;
      end
    end else begin
      spriteYRegs_26 <= _GEN_39;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_27 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_27 <= _GEN_41;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_27 <= _GEN_300;
      end else begin
        spriteYRegs_27 <= _GEN_41;
      end
    end else begin
      spriteYRegs_27 <= _GEN_41;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_28 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_28 <= _GEN_43;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_28 <= _GEN_305;
      end else begin
        spriteYRegs_28 <= _GEN_43;
      end
    end else begin
      spriteYRegs_28 <= _GEN_43;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_29 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_29 <= _GEN_45;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_29 <= _GEN_310;
      end else begin
        spriteYRegs_29 <= _GEN_45;
      end
    end else begin
      spriteYRegs_29 <= _GEN_45;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_30 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_30 <= _GEN_47;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_30 <= _GEN_315;
      end else begin
        spriteYRegs_30 <= _GEN_47;
      end
    end else begin
      spriteYRegs_30 <= _GEN_47;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_31 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_31 <= _GEN_49;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_31 <= _GEN_320;
      end else begin
        spriteYRegs_31 <= _GEN_49;
      end
    end else begin
      spriteYRegs_31 <= _GEN_49;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_32 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_32 <= _GEN_51;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_32 <= _GEN_325;
      end else begin
        spriteYRegs_32 <= _GEN_51;
      end
    end else begin
      spriteYRegs_32 <= _GEN_51;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_33 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_33 <= _GEN_53;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_33 <= _GEN_330;
      end else begin
        spriteYRegs_33 <= _GEN_53;
      end
    end else begin
      spriteYRegs_33 <= _GEN_53;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_34 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_34 <= _GEN_55;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_34 <= _GEN_335;
      end else begin
        spriteYRegs_34 <= _GEN_55;
      end
    end else begin
      spriteYRegs_34 <= _GEN_55;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_35 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_35 <= _GEN_57;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_35 <= _GEN_340;
      end else begin
        spriteYRegs_35 <= _GEN_57;
      end
    end else begin
      spriteYRegs_35 <= _GEN_57;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_36 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_36 <= _GEN_59;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_36 <= _GEN_345;
      end else begin
        spriteYRegs_36 <= _GEN_59;
      end
    end else begin
      spriteYRegs_36 <= _GEN_59;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_37 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_37 <= _GEN_61;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_37 <= _GEN_350;
      end else begin
        spriteYRegs_37 <= _GEN_61;
      end
    end else begin
      spriteYRegs_37 <= _GEN_61;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_38 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_38 <= _GEN_63;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_38 <= _GEN_355;
      end else begin
        spriteYRegs_38 <= _GEN_63;
      end
    end else begin
      spriteYRegs_38 <= _GEN_63;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_39 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_39 <= _GEN_65;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_39 <= _GEN_360;
      end else begin
        spriteYRegs_39 <= _GEN_65;
      end
    end else begin
      spriteYRegs_39 <= _GEN_65;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_40 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_40 <= _GEN_67;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_40 <= _GEN_365;
      end else begin
        spriteYRegs_40 <= _GEN_67;
      end
    end else begin
      spriteYRegs_40 <= _GEN_67;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_41 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_41 <= _GEN_69;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_41 <= _GEN_370;
      end else begin
        spriteYRegs_41 <= _GEN_69;
      end
    end else begin
      spriteYRegs_41 <= _GEN_69;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_42 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_42 <= _GEN_71;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_42 <= _GEN_375;
      end else begin
        spriteYRegs_42 <= _GEN_71;
      end
    end else begin
      spriteYRegs_42 <= _GEN_71;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_43 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_43 <= _GEN_73;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_43 <= _GEN_380;
      end else begin
        spriteYRegs_43 <= _GEN_73;
      end
    end else begin
      spriteYRegs_43 <= _GEN_73;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_44 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_44 <= _GEN_75;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_44 <= _GEN_385;
      end else begin
        spriteYRegs_44 <= _GEN_75;
      end
    end else begin
      spriteYRegs_44 <= _GEN_75;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_45 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_45 <= _GEN_77;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        spriteYRegs_45 <= _GEN_390;
      end else begin
        spriteYRegs_45 <= _GEN_77;
      end
    end else begin
      spriteYRegs_45 <= _GEN_77;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_46 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_46 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_47 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_47 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_48 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_48 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_49 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_49 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_50 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_50 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_51 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_51 <= 10'shc8; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_52 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_52 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_53 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_53 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_54 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_54 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_55 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_55 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_56 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_56 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_57 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_57 <= 10'sh104; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_58 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_58 <= _GEN_103;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 594:29]
        spriteYRegs_58 <= spriteYRegs_58_REG; // @[\\src\\main\\scala\\GameLogic.scala 596:25]
      end else begin
        spriteYRegs_58 <= _GEN_1244;
      end
    end else begin
      spriteYRegs_58 <= _GEN_103;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_59 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_59 <= _GEN_105;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 594:29]
        spriteYRegs_59 <= spriteYRegs_59_REG; // @[\\src\\main\\scala\\GameLogic.scala 598:25]
      end else begin
        spriteYRegs_59 <= _GEN_1245;
      end
    end else begin
      spriteYRegs_59 <= _GEN_105;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_60 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteYRegs_60 <= _GEN_107;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 594:29]
        spriteYRegs_60 <= spriteYRegs_60_REG; // @[\\src\\main\\scala\\GameLogic.scala 600:25]
      end else begin
        spriteYRegs_60 <= _GEN_1246;
      end
    end else begin
      spriteYRegs_60 <= _GEN_107;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_61 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_61 <= 10'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_62 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_62 <= 10'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 122:28]
      spriteYRegs_63 <= 10'sh0; // @[\\src\\main\\scala\\GameLogic.scala 122:28]
    end else if (initializePositions) begin // @[\\src\\main\\scala\\GameLogic.scala 131:29]
      spriteYRegs_63 <= 10'sh14; // @[\\src\\main\\scala\\GameLogic.scala 162:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_3 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        spriteVisibleRegs_3 <= _GEN_139;
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_3 <= _GEN_601;
      end else begin
        spriteVisibleRegs_3 <= _GEN_995;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_3 <= _GEN_1285;
    end else begin
      spriteVisibleRegs_3 <= _GEN_1369;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_4 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_4 <= _GEN_602;
        end else begin
          spriteVisibleRegs_4 <= _GEN_996;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_5 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_5 <= _GEN_603;
        end else begin
          spriteVisibleRegs_5 <= _GEN_997;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_6 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_6 <= _GEN_604;
        end else begin
          spriteVisibleRegs_6 <= _GEN_998;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_7 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_7 <= _GEN_605;
        end else begin
          spriteVisibleRegs_7 <= _GEN_999;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        spriteVisibleRegs_7 <= _GEN_1286;
      end else begin
        spriteVisibleRegs_7 <= _GEN_1370;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_8 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_8 <= _GEN_606;
        end else begin
          spriteVisibleRegs_8 <= _GEN_1000;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        spriteVisibleRegs_8 <= _GEN_1287;
      end else begin
        spriteVisibleRegs_8 <= _GEN_1371;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_9 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_9 <= _GEN_607;
        end else begin
          spriteVisibleRegs_9 <= _GEN_1001;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        spriteVisibleRegs_9 <= _GEN_1288;
      end else begin
        spriteVisibleRegs_9 <= _GEN_1372;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_10 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_10 <= _GEN_608;
        end else begin
          spriteVisibleRegs_10 <= _GEN_1002;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        spriteVisibleRegs_10 <= _GEN_1289;
      end else begin
        spriteVisibleRegs_10 <= _GEN_1373;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_11 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_11 <= _GEN_609;
        end else begin
          spriteVisibleRegs_11 <= _GEN_1003;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        spriteVisibleRegs_11 <= _GEN_1290;
      end else begin
        spriteVisibleRegs_11 <= _GEN_1374;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_12 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_12 <= _GEN_610;
        end else begin
          spriteVisibleRegs_12 <= _GEN_1004;
        end
      end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        spriteVisibleRegs_12 <= _GEN_1291;
      end else begin
        spriteVisibleRegs_12 <= _GEN_1375;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_13 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T_792) begin // @[\\src\\main\\scala\\GameLogic.scala 540:9]
          spriteVisibleRegs_13 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 541:31]
        end else begin
          spriteVisibleRegs_13 <= _GEN_1071;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_14 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_14 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 297:27]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 555:24]
        spriteVisibleRegs_14 <= _GEN_1170;
      end else begin
        spriteVisibleRegs_14 <= _GEN_1072;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_14 <= _GEN_1376;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_15 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
          spriteVisibleRegs_15 <= _GEN_613;
        end else begin
          spriteVisibleRegs_15 <= _GEN_1007;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_16 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_16 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_16 <= _GEN_614;
      end else begin
        spriteVisibleRegs_16 <= _GEN_1008;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_17 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_17 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_17 <= _GEN_615;
      end else begin
        spriteVisibleRegs_17 <= _GEN_1009;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_18 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_18 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_18 <= _GEN_616;
      end else begin
        spriteVisibleRegs_18 <= _GEN_1010;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_19 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_19 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_19 <= _GEN_617;
      end else begin
        spriteVisibleRegs_19 <= _GEN_1011;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_20 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_20 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_20 <= _GEN_618;
      end else begin
        spriteVisibleRegs_20 <= _GEN_1012;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_21 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_21 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_21 <= _GEN_619;
      end else begin
        spriteVisibleRegs_21 <= _GEN_1013;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_22 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_22 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_22 <= _GEN_620;
      end else begin
        spriteVisibleRegs_22 <= _GEN_1014;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_23 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_23 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_23 <= _GEN_621;
      end else begin
        spriteVisibleRegs_23 <= _GEN_1015;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_24 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_24 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_24 <= _GEN_622;
      end else begin
        spriteVisibleRegs_24 <= _GEN_1016;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_25 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_25 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_25 <= _GEN_623;
      end else begin
        spriteVisibleRegs_25 <= _GEN_1017;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_26 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_26 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_26 <= _GEN_624;
      end else begin
        spriteVisibleRegs_26 <= _GEN_1018;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_27 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_27 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_27 <= _GEN_625;
      end else begin
        spriteVisibleRegs_27 <= _GEN_1019;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_28 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_28 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_28 <= _GEN_626;
      end else begin
        spriteVisibleRegs_28 <= _GEN_1020;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_29 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_29 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_29 <= _GEN_627;
      end else begin
        spriteVisibleRegs_29 <= _GEN_1021;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_30 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_30 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_30 <= _GEN_628;
      end else begin
        spriteVisibleRegs_30 <= _GEN_1022;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_31 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_31 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_31 <= _GEN_629;
      end else begin
        spriteVisibleRegs_31 <= _GEN_1023;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_32 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_32 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_32 <= _GEN_630;
      end else begin
        spriteVisibleRegs_32 <= _GEN_1024;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_33 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_33 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_33 <= _GEN_631;
      end else begin
        spriteVisibleRegs_33 <= _GEN_1025;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_34 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_34 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_34 <= _GEN_632;
      end else begin
        spriteVisibleRegs_34 <= _GEN_1026;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_35 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_35 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_35 <= _GEN_633;
      end else begin
        spriteVisibleRegs_35 <= _GEN_1027;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_36 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_36 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_36 <= _GEN_634;
      end else begin
        spriteVisibleRegs_36 <= _GEN_1028;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_37 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_37 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_37 <= _GEN_635;
      end else begin
        spriteVisibleRegs_37 <= _GEN_1029;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_38 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_38 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_38 <= _GEN_636;
      end else begin
        spriteVisibleRegs_38 <= _GEN_1030;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_39 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_39 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_39 <= _GEN_637;
      end else begin
        spriteVisibleRegs_39 <= _GEN_1031;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_40 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_40 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_40 <= _GEN_638;
      end else begin
        spriteVisibleRegs_40 <= _GEN_1032;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_41 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_41 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_41 <= _GEN_639;
      end else begin
        spriteVisibleRegs_41 <= _GEN_1033;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_42 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_42 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_42 <= _GEN_640;
      end else begin
        spriteVisibleRegs_42 <= _GEN_1034;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_43 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_43 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_43 <= _GEN_641;
      end else begin
        spriteVisibleRegs_43 <= _GEN_1035;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_44 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_44 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_44 <= _GEN_642;
      end else begin
        spriteVisibleRegs_44 <= _GEN_1036;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_45 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_45 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 301:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_45 <= _GEN_643;
      end else begin
        spriteVisibleRegs_45 <= _GEN_1037;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_46 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_46 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_46 <= _GEN_644;
      end else begin
        spriteVisibleRegs_46 <= _GEN_1038;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_46 <= _GEN_1385;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_47 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_47 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_47 <= _GEN_645;
      end else begin
        spriteVisibleRegs_47 <= _GEN_1039;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_47 <= _GEN_1386;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_48 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_48 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_48 <= _GEN_646;
      end else begin
        spriteVisibleRegs_48 <= _GEN_1040;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_48 <= _GEN_1387;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_49 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_49 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_49 <= _GEN_647;
      end else begin
        spriteVisibleRegs_49 <= _GEN_1041;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_49 <= _GEN_1388;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_50 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_50 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_50 <= _GEN_648;
      end else begin
        spriteVisibleRegs_50 <= _GEN_1042;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_50 <= _GEN_1389;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_51 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_51 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_51 <= _GEN_649;
      end else begin
        spriteVisibleRegs_51 <= _GEN_1043;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_51 <= _GEN_1390;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_52 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_52 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_52 <= _GEN_650;
      end else begin
        spriteVisibleRegs_52 <= _GEN_1044;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_52 <= _GEN_1391;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_53 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_53 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_53 <= _GEN_651;
      end else begin
        spriteVisibleRegs_53 <= _GEN_1045;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_53 <= _GEN_1392;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_54 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_54 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_54 <= _GEN_652;
      end else begin
        spriteVisibleRegs_54 <= _GEN_1046;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_54 <= _GEN_1393;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_55 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_55 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_55 <= _GEN_653;
      end else begin
        spriteVisibleRegs_55 <= _GEN_1047;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_55 <= _GEN_1394;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_56 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_56 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_56 <= _GEN_654;
      end else begin
        spriteVisibleRegs_56 <= _GEN_1048;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_56 <= _GEN_1395;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_57 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spriteVisibleRegs_57 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 306:28]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_57 <= _GEN_655;
      end else begin
        spriteVisibleRegs_57 <= _GEN_1049;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_57 <= _GEN_1396;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_58 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        spriteVisibleRegs_58 <= _T_83;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_59 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        spriteVisibleRegs_59 <= _T_83;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_60 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        spriteVisibleRegs_60 <= _T_83;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_61 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_61 <= _GEN_123;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_61 <= _GEN_659;
      end else begin
        spriteVisibleRegs_61 <= _GEN_1053;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_61 <= _GEN_123;
    end else begin
      spriteVisibleRegs_61 <= _GEN_1377;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_62 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_62 <= _GEN_124;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_62 <= _GEN_660;
      end else begin
        spriteVisibleRegs_62 <= _GEN_1054;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_62 <= _GEN_124;
    end else begin
      spriteVisibleRegs_62 <= _GEN_1378;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 125:34]
      spriteVisibleRegs_63 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 125:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_63 <= _GEN_125;
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spriteVisibleRegs_63 <= _GEN_661;
      end else begin
        spriteVisibleRegs_63 <= _GEN_1055;
      end
    end else if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spriteVisibleRegs_63 <= _GEN_125;
    end else begin
      spriteVisibleRegs_63 <= _GEN_1379;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_0 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_0 <= _GEN_346;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_1 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_1 <= _GEN_351;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_2 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_2 <= _GEN_356;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_3 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_3 <= _GEN_361;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_4 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_4 <= _GEN_366;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_5 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_5 <= _GEN_371;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_6 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_6 <= _GEN_376;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_7 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_7 <= _GEN_381;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_8 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_8 <= _GEN_386;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 126:36]
      spriteScaleTypeRegs_9 <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 126:36]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
          spriteScaleTypeRegs_9 <= _GEN_391;
        end
      end
    end
    initializePositions <= reset | _GEN_1674; // @[\\src\\main\\scala\\GameLogic.scala 130:{36,36}]
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 168:42]
      sprite58ScaleUpHorizontal <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 168:42]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        sprite58ScaleUpHorizontal <= _GEN_1254;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 169:40]
      sprite58ScaleUpVertical <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 169:40]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        sprite58ScaleUpVertical <= _GEN_1257;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 170:42]
      sprite59ScaleUpHorizontal <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 170:42]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        sprite59ScaleUpHorizontal <= _GEN_1255;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 171:40]
      sprite59ScaleUpVertical <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 171:40]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        sprite59ScaleUpVertical <= _GEN_1258;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 172:42]
      sprite60ScaleUpHorizontal <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 172:42]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        sprite60ScaleUpHorizontal <= _GEN_1256;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 173:40]
      sprite60ScaleUpVertical <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 173:40]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        sprite60ScaleUpVertical <= _GEN_1259;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 201:28]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 201:28]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
          viewBoxXReg <= _GEN_1380;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 202:28]
      viewBoxYReg <= 9'h0; // @[\\src\\main\\scala\\GameLogic.scala 202:28]
    end else if (!(3'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
          viewBoxYReg <= _GEN_1381;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 211:23]
      lvlReg <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 211:23]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          lvlReg <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 282:12]
        end
      end
    end else if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (3'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        lvlReg <= _GEN_1292;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 222:25]
      livesReg <= 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 222:25]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          livesReg <= 3'h3; // @[\\src\\main\\scala\\GameLogic.scala 283:14]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 555:24]
        livesReg <= _GEN_1171;
      end else begin
        livesReg <= _GEN_1159;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 225:29]
      extraLifeCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 225:29]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          extraLifeCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 287:18]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (_T) begin // @[\\src\\main\\scala\\GameLogic.scala 359:29]
        extraLifeCnt <= _GEN_396;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 231:34]
      spawnDelayCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 231:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          spawnDelayCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 285:23]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        spawnDelayCounter <= _GEN_663;
      end else begin
        spawnDelayCounter <= _GEN_1057;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      spawnDelayCounter <= _GEN_1366;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 232:34]
      nextSpriteToSpawn <= 6'h0; // @[\\src\\main\\scala\\GameLogic.scala 232:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          nextSpriteToSpawn <= 6'h0; // @[\\src\\main\\scala\\GameLogic.scala 286:23]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (lvlReg == 2'h1) begin // @[\\src\\main\\scala\\GameLogic.scala 450:28]
        nextSpriteToSpawn <= _GEN_662;
      end else begin
        nextSpriteToSpawn <= _GEN_1056;
      end
    end else if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      nextSpriteToSpawn <= _GEN_1365;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 235:24]
      starCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 235:24]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          starCnt <= 10'h0; // @[\\src\\main\\scala\\GameLogic.scala 288:13]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (starCnt == 10'h0) begin // @[\\src\\main\\scala\\GameLogic.scala 594:29]
        starCnt <= _starCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 607:17]
      end else begin
        starCnt <= _GEN_1247;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 238:34]
      collisionDetected <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 238:34]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          collisionDetected <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 289:23]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 555:24]
        collisionDetected <= _GEN_1173;
      end else begin
        collisionDetected <= _GEN_1156;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 239:29]
      blinkCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 239:29]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          blinkCounter <= 8'h0; // @[\\src\\main\\scala\\GameLogic.scala 291:18]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 555:24]
        blinkCounter <= _GEN_1165;
      end else begin
        blinkCounter <= _GEN_1161;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 240:27]
      blinkTimes <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 240:27]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          blinkTimes <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 292:16]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 555:24]
        blinkTimes <= _GEN_1166;
      end else begin
        blinkTimes <= _GEN_1162;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 241:27]
      isBlinking <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 241:27]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          isBlinking <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 290:16]
        end
      end
    end else if (3'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (isBlinking) begin // @[\\src\\main\\scala\\GameLogic.scala 555:24]
        isBlinking <= _GEN_1169;
      end else begin
        isBlinking <= _GEN_1160;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 247:38]
      gameOverReturnPressed <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 247:38]
    end else if (3'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (io_newFrame) begin // @[\\src\\main\\scala\\GameLogic.scala 338:25]
        if (gameOverReturnPressed) begin // @[\\src\\main\\scala\\GameLogic.scala 339:37]
          gameOverReturnPressed <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 341:33]
        end
      end
    end else if (!(3'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
      if (!(3'h2 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 336:20]
        gameOverReturnPressed <= _GEN_1397;
      end
    end
    spriteXRegs_58_REG <= $signed(spriteXRegs_59) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 595:52]
    spriteYRegs_58_REG <= $signed(spriteYRegs_59) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 596:52]
    spriteXRegs_59_REG <= $signed(spriteXRegs_60) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 597:52]
    spriteYRegs_59_REG <= $signed(spriteYRegs_60) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 598:52]
    spriteXRegs_60_REG <= $signed(spriteXRegs_58) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 599:52]
    spriteYRegs_60_REG <= $signed(spriteYRegs_58) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 600:52]
    spriteXRegs_58_REG_1 <= $signed(spriteXRegs_59) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 623:52]
    spriteYRegs_58_REG_1 <= $signed(spriteYRegs_59) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 624:52]
    spriteXRegs_59_REG_1 <= $signed(spriteXRegs_60) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 625:52]
    spriteYRegs_59_REG_1 <= $signed(spriteYRegs_60) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 626:52]
    spriteXRegs_60_REG_1 <= $signed(spriteXRegs_58) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 627:52]
    spriteYRegs_60_REG_1 <= $signed(spriteYRegs_58) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 628:52]
    spriteXRegs_58_REG_2 <= $signed(spriteXRegs_59) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 651:52]
    spriteYRegs_58_REG_2 <= $signed(spriteYRegs_59) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 652:52]
    spriteXRegs_59_REG_2 <= $signed(spriteXRegs_60) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 653:52]
    spriteYRegs_59_REG_2 <= $signed(spriteYRegs_60) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 654:52]
    spriteXRegs_60_REG_2 <= $signed(spriteXRegs_58) - 11'sh10; // @[\\src\\main\\scala\\GameLogic.scala 655:52]
    spriteYRegs_60_REG_2 <= $signed(spriteYRegs_58) - 10'sh10; // @[\\src\\main\\scala\\GameLogic.scala 656:52]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  spriteXRegs_3 = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  spriteXRegs_7 = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  spriteXRegs_8 = _RAND_3[10:0];
  _RAND_4 = {1{`RANDOM}};
  spriteXRegs_9 = _RAND_4[10:0];
  _RAND_5 = {1{`RANDOM}};
  spriteXRegs_10 = _RAND_5[10:0];
  _RAND_6 = {1{`RANDOM}};
  spriteXRegs_11 = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  spriteXRegs_12 = _RAND_7[10:0];
  _RAND_8 = {1{`RANDOM}};
  spriteXRegs_13 = _RAND_8[10:0];
  _RAND_9 = {1{`RANDOM}};
  spriteXRegs_14 = _RAND_9[10:0];
  _RAND_10 = {1{`RANDOM}};
  spriteXRegs_16 = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  spriteXRegs_17 = _RAND_11[10:0];
  _RAND_12 = {1{`RANDOM}};
  spriteXRegs_18 = _RAND_12[10:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXRegs_19 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXRegs_20 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXRegs_21 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXRegs_22 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXRegs_23 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXRegs_24 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXRegs_25 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteXRegs_26 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  spriteXRegs_27 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  spriteXRegs_28 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  spriteXRegs_29 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  spriteXRegs_30 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  spriteXRegs_31 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  spriteXRegs_32 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  spriteXRegs_33 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  spriteXRegs_34 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  spriteXRegs_35 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  spriteXRegs_36 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  spriteXRegs_37 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  spriteXRegs_38 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  spriteXRegs_39 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  spriteXRegs_40 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  spriteXRegs_41 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  spriteXRegs_42 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  spriteXRegs_43 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  spriteXRegs_44 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  spriteXRegs_45 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  spriteXRegs_46 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  spriteXRegs_47 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  spriteXRegs_48 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  spriteXRegs_49 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  spriteXRegs_50 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  spriteXRegs_51 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  spriteXRegs_52 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  spriteXRegs_53 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  spriteXRegs_54 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  spriteXRegs_55 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  spriteXRegs_56 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  spriteXRegs_57 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  spriteXRegs_58 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  spriteXRegs_59 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  spriteXRegs_60 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  spriteXRegs_61 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  spriteXRegs_62 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  spriteXRegs_63 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  spriteYRegs_3 = _RAND_58[9:0];
  _RAND_59 = {1{`RANDOM}};
  spriteYRegs_7 = _RAND_59[9:0];
  _RAND_60 = {1{`RANDOM}};
  spriteYRegs_8 = _RAND_60[9:0];
  _RAND_61 = {1{`RANDOM}};
  spriteYRegs_9 = _RAND_61[9:0];
  _RAND_62 = {1{`RANDOM}};
  spriteYRegs_10 = _RAND_62[9:0];
  _RAND_63 = {1{`RANDOM}};
  spriteYRegs_11 = _RAND_63[9:0];
  _RAND_64 = {1{`RANDOM}};
  spriteYRegs_12 = _RAND_64[9:0];
  _RAND_65 = {1{`RANDOM}};
  spriteYRegs_13 = _RAND_65[9:0];
  _RAND_66 = {1{`RANDOM}};
  spriteYRegs_14 = _RAND_66[9:0];
  _RAND_67 = {1{`RANDOM}};
  spriteYRegs_16 = _RAND_67[9:0];
  _RAND_68 = {1{`RANDOM}};
  spriteYRegs_17 = _RAND_68[9:0];
  _RAND_69 = {1{`RANDOM}};
  spriteYRegs_18 = _RAND_69[9:0];
  _RAND_70 = {1{`RANDOM}};
  spriteYRegs_19 = _RAND_70[9:0];
  _RAND_71 = {1{`RANDOM}};
  spriteYRegs_20 = _RAND_71[9:0];
  _RAND_72 = {1{`RANDOM}};
  spriteYRegs_21 = _RAND_72[9:0];
  _RAND_73 = {1{`RANDOM}};
  spriteYRegs_22 = _RAND_73[9:0];
  _RAND_74 = {1{`RANDOM}};
  spriteYRegs_23 = _RAND_74[9:0];
  _RAND_75 = {1{`RANDOM}};
  spriteYRegs_24 = _RAND_75[9:0];
  _RAND_76 = {1{`RANDOM}};
  spriteYRegs_25 = _RAND_76[9:0];
  _RAND_77 = {1{`RANDOM}};
  spriteYRegs_26 = _RAND_77[9:0];
  _RAND_78 = {1{`RANDOM}};
  spriteYRegs_27 = _RAND_78[9:0];
  _RAND_79 = {1{`RANDOM}};
  spriteYRegs_28 = _RAND_79[9:0];
  _RAND_80 = {1{`RANDOM}};
  spriteYRegs_29 = _RAND_80[9:0];
  _RAND_81 = {1{`RANDOM}};
  spriteYRegs_30 = _RAND_81[9:0];
  _RAND_82 = {1{`RANDOM}};
  spriteYRegs_31 = _RAND_82[9:0];
  _RAND_83 = {1{`RANDOM}};
  spriteYRegs_32 = _RAND_83[9:0];
  _RAND_84 = {1{`RANDOM}};
  spriteYRegs_33 = _RAND_84[9:0];
  _RAND_85 = {1{`RANDOM}};
  spriteYRegs_34 = _RAND_85[9:0];
  _RAND_86 = {1{`RANDOM}};
  spriteYRegs_35 = _RAND_86[9:0];
  _RAND_87 = {1{`RANDOM}};
  spriteYRegs_36 = _RAND_87[9:0];
  _RAND_88 = {1{`RANDOM}};
  spriteYRegs_37 = _RAND_88[9:0];
  _RAND_89 = {1{`RANDOM}};
  spriteYRegs_38 = _RAND_89[9:0];
  _RAND_90 = {1{`RANDOM}};
  spriteYRegs_39 = _RAND_90[9:0];
  _RAND_91 = {1{`RANDOM}};
  spriteYRegs_40 = _RAND_91[9:0];
  _RAND_92 = {1{`RANDOM}};
  spriteYRegs_41 = _RAND_92[9:0];
  _RAND_93 = {1{`RANDOM}};
  spriteYRegs_42 = _RAND_93[9:0];
  _RAND_94 = {1{`RANDOM}};
  spriteYRegs_43 = _RAND_94[9:0];
  _RAND_95 = {1{`RANDOM}};
  spriteYRegs_44 = _RAND_95[9:0];
  _RAND_96 = {1{`RANDOM}};
  spriteYRegs_45 = _RAND_96[9:0];
  _RAND_97 = {1{`RANDOM}};
  spriteYRegs_46 = _RAND_97[9:0];
  _RAND_98 = {1{`RANDOM}};
  spriteYRegs_47 = _RAND_98[9:0];
  _RAND_99 = {1{`RANDOM}};
  spriteYRegs_48 = _RAND_99[9:0];
  _RAND_100 = {1{`RANDOM}};
  spriteYRegs_49 = _RAND_100[9:0];
  _RAND_101 = {1{`RANDOM}};
  spriteYRegs_50 = _RAND_101[9:0];
  _RAND_102 = {1{`RANDOM}};
  spriteYRegs_51 = _RAND_102[9:0];
  _RAND_103 = {1{`RANDOM}};
  spriteYRegs_52 = _RAND_103[9:0];
  _RAND_104 = {1{`RANDOM}};
  spriteYRegs_53 = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  spriteYRegs_54 = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  spriteYRegs_55 = _RAND_106[9:0];
  _RAND_107 = {1{`RANDOM}};
  spriteYRegs_56 = _RAND_107[9:0];
  _RAND_108 = {1{`RANDOM}};
  spriteYRegs_57 = _RAND_108[9:0];
  _RAND_109 = {1{`RANDOM}};
  spriteYRegs_58 = _RAND_109[9:0];
  _RAND_110 = {1{`RANDOM}};
  spriteYRegs_59 = _RAND_110[9:0];
  _RAND_111 = {1{`RANDOM}};
  spriteYRegs_60 = _RAND_111[9:0];
  _RAND_112 = {1{`RANDOM}};
  spriteYRegs_61 = _RAND_112[9:0];
  _RAND_113 = {1{`RANDOM}};
  spriteYRegs_62 = _RAND_113[9:0];
  _RAND_114 = {1{`RANDOM}};
  spriteYRegs_63 = _RAND_114[9:0];
  _RAND_115 = {1{`RANDOM}};
  spriteVisibleRegs_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  spriteVisibleRegs_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  spriteVisibleRegs_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  spriteVisibleRegs_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  spriteVisibleRegs_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  spriteVisibleRegs_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  spriteVisibleRegs_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  spriteVisibleRegs_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  spriteVisibleRegs_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  spriteVisibleRegs_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  spriteVisibleRegs_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  spriteVisibleRegs_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  spriteVisibleRegs_15 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  spriteVisibleRegs_16 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  spriteVisibleRegs_17 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  spriteVisibleRegs_18 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  spriteVisibleRegs_19 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  spriteVisibleRegs_20 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  spriteVisibleRegs_21 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  spriteVisibleRegs_22 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  spriteVisibleRegs_23 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  spriteVisibleRegs_24 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  spriteVisibleRegs_25 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  spriteVisibleRegs_26 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  spriteVisibleRegs_27 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  spriteVisibleRegs_28 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  spriteVisibleRegs_29 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  spriteVisibleRegs_30 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  spriteVisibleRegs_31 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  spriteVisibleRegs_32 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  spriteVisibleRegs_33 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  spriteVisibleRegs_34 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  spriteVisibleRegs_35 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  spriteVisibleRegs_36 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  spriteVisibleRegs_37 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  spriteVisibleRegs_38 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  spriteVisibleRegs_39 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  spriteVisibleRegs_40 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  spriteVisibleRegs_41 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  spriteVisibleRegs_42 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  spriteVisibleRegs_43 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  spriteVisibleRegs_44 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  spriteVisibleRegs_45 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  spriteVisibleRegs_46 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  spriteVisibleRegs_47 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  spriteVisibleRegs_48 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  spriteVisibleRegs_49 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  spriteVisibleRegs_50 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  spriteVisibleRegs_51 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  spriteVisibleRegs_52 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  spriteVisibleRegs_53 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  spriteVisibleRegs_54 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  spriteVisibleRegs_55 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  spriteVisibleRegs_56 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  spriteVisibleRegs_57 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  spriteVisibleRegs_58 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  spriteVisibleRegs_59 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  spriteVisibleRegs_60 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  spriteVisibleRegs_61 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  spriteVisibleRegs_62 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  spriteVisibleRegs_63 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  spriteScaleTypeRegs_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  spriteScaleTypeRegs_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  spriteScaleTypeRegs_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  spriteScaleTypeRegs_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  spriteScaleTypeRegs_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  spriteScaleTypeRegs_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  spriteScaleTypeRegs_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  spriteScaleTypeRegs_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  spriteScaleTypeRegs_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  spriteScaleTypeRegs_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  initializePositions = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  sprite58ScaleUpHorizontal = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  sprite58ScaleUpVertical = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  sprite59ScaleUpHorizontal = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  sprite59ScaleUpVertical = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  sprite60ScaleUpHorizontal = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  sprite60ScaleUpVertical = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  viewBoxXReg = _RAND_193[9:0];
  _RAND_194 = {1{`RANDOM}};
  viewBoxYReg = _RAND_194[8:0];
  _RAND_195 = {1{`RANDOM}};
  lvlReg = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  livesReg = _RAND_196[2:0];
  _RAND_197 = {1{`RANDOM}};
  extraLifeCnt = _RAND_197[9:0];
  _RAND_198 = {1{`RANDOM}};
  spawnDelayCounter = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  nextSpriteToSpawn = _RAND_199[5:0];
  _RAND_200 = {1{`RANDOM}};
  starCnt = _RAND_200[9:0];
  _RAND_201 = {1{`RANDOM}};
  collisionDetected = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  blinkCounter = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  blinkTimes = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  isBlinking = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  gameOverReturnPressed = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  spriteXRegs_58_REG = _RAND_206[10:0];
  _RAND_207 = {1{`RANDOM}};
  spriteYRegs_58_REG = _RAND_207[9:0];
  _RAND_208 = {1{`RANDOM}};
  spriteXRegs_59_REG = _RAND_208[10:0];
  _RAND_209 = {1{`RANDOM}};
  spriteYRegs_59_REG = _RAND_209[9:0];
  _RAND_210 = {1{`RANDOM}};
  spriteXRegs_60_REG = _RAND_210[10:0];
  _RAND_211 = {1{`RANDOM}};
  spriteYRegs_60_REG = _RAND_211[9:0];
  _RAND_212 = {1{`RANDOM}};
  spriteXRegs_58_REG_1 = _RAND_212[10:0];
  _RAND_213 = {1{`RANDOM}};
  spriteYRegs_58_REG_1 = _RAND_213[9:0];
  _RAND_214 = {1{`RANDOM}};
  spriteXRegs_59_REG_1 = _RAND_214[10:0];
  _RAND_215 = {1{`RANDOM}};
  spriteYRegs_59_REG_1 = _RAND_215[9:0];
  _RAND_216 = {1{`RANDOM}};
  spriteXRegs_60_REG_1 = _RAND_216[10:0];
  _RAND_217 = {1{`RANDOM}};
  spriteYRegs_60_REG_1 = _RAND_217[9:0];
  _RAND_218 = {1{`RANDOM}};
  spriteXRegs_58_REG_2 = _RAND_218[10:0];
  _RAND_219 = {1{`RANDOM}};
  spriteYRegs_58_REG_2 = _RAND_219[9:0];
  _RAND_220 = {1{`RANDOM}};
  spriteXRegs_59_REG_2 = _RAND_220[10:0];
  _RAND_221 = {1{`RANDOM}};
  spriteYRegs_59_REG_2 = _RAND_221[9:0];
  _RAND_222 = {1{`RANDOM}};
  spriteXRegs_60_REG_2 = _RAND_222[10:0];
  _RAND_223 = {1{`RANDOM}};
  spriteYRegs_60_REG_2 = _RAND_223[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GameTop(
  input        clock,
  input        reset,
  input        io_btnC, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnU, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnL, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnR, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnD, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaRed, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaBlue, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaGreen, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_Hsync, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_Vsync, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_missingFrameError, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_viewBoxOutOfRangeError // @[\\src\\main\\scala\\GameTop.scala 14:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  graphicEngineVGA_clock; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_reset; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_46; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_47; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_48; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_49; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_50; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_51; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_52; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_53; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_54; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_55; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_56; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_57; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_61; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_62; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_63; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_46; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_47; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_48; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_49; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_50; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_51; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_52; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_53; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_54; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_55; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_56; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_57; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_61; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_62; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_63; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_46; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_47; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_48; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_49; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_50; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_51; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_52; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_53; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_54; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_55; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_56; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_57; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_61; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_62; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_63; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [8:0] graphicEngineVGA_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_missingFrameError; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaRed; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaBlue; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaGreen; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Hsync; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Vsync; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  soundEngine_clock; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  soundEngine_reset; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  gameLogic_clock; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_reset; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnC; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnU; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnL; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnR; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnD; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_46; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_47; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_48; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_49; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_50; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_51; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_52; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_53; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_54; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_55; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_56; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_57; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_61; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_62; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_63; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_46; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_47; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_48; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_49; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_50; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_51; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_52; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_53; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_54; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_55; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_56; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_57; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_61; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_62; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_63; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_46; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_47; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_48; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_49; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_50; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_51; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_52; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_53; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_54; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_55; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_56; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_57; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_61; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_62; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_63; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [8:0] gameLogic_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  reg [20:0] debounceCounter; // @[\\src\\main\\scala\\GameTop.scala 68:32]
  wire  debounceSampleEn = debounceCounter == 21'h1e847f; // @[\\src\\main\\scala\\GameTop.scala 70:24]
  wire [20:0] _debounceCounter_T_1 = debounceCounter + 21'h1; // @[\\src\\main\\scala\\GameTop.scala 74:40]
  reg [21:0] resetReleaseCounter; // @[\\src\\main\\scala\\GameTop.scala 81:36]
  wire [21:0] _resetReleaseCounter_T_1 = resetReleaseCounter + 22'h1; // @[\\src\\main\\scala\\GameTop.scala 87:48]
  reg  btnCState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnCState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnCState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnCState; // @[\\src\\main\\scala\\GameTop.scala 93:28]
  reg  btnUState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState; // @[\\src\\main\\scala\\GameTop.scala 94:28]
  reg  btnLState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState; // @[\\src\\main\\scala\\GameTop.scala 95:28]
  reg  btnRState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState; // @[\\src\\main\\scala\\GameTop.scala 96:28]
  reg  btnDState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState; // @[\\src\\main\\scala\\GameTop.scala 97:28]
  GraphicEngineVGA graphicEngineVGA ( // @[\\src\\main\\scala\\GameTop.scala 46:32]
    .clock(graphicEngineVGA_clock),
    .reset(graphicEngineVGA_reset),
    .io_spriteXPosition_3(graphicEngineVGA_io_spriteXPosition_3),
    .io_spriteXPosition_7(graphicEngineVGA_io_spriteXPosition_7),
    .io_spriteXPosition_8(graphicEngineVGA_io_spriteXPosition_8),
    .io_spriteXPosition_9(graphicEngineVGA_io_spriteXPosition_9),
    .io_spriteXPosition_10(graphicEngineVGA_io_spriteXPosition_10),
    .io_spriteXPosition_11(graphicEngineVGA_io_spriteXPosition_11),
    .io_spriteXPosition_12(graphicEngineVGA_io_spriteXPosition_12),
    .io_spriteXPosition_13(graphicEngineVGA_io_spriteXPosition_13),
    .io_spriteXPosition_14(graphicEngineVGA_io_spriteXPosition_14),
    .io_spriteXPosition_16(graphicEngineVGA_io_spriteXPosition_16),
    .io_spriteXPosition_17(graphicEngineVGA_io_spriteXPosition_17),
    .io_spriteXPosition_18(graphicEngineVGA_io_spriteXPosition_18),
    .io_spriteXPosition_19(graphicEngineVGA_io_spriteXPosition_19),
    .io_spriteXPosition_20(graphicEngineVGA_io_spriteXPosition_20),
    .io_spriteXPosition_21(graphicEngineVGA_io_spriteXPosition_21),
    .io_spriteXPosition_22(graphicEngineVGA_io_spriteXPosition_22),
    .io_spriteXPosition_23(graphicEngineVGA_io_spriteXPosition_23),
    .io_spriteXPosition_24(graphicEngineVGA_io_spriteXPosition_24),
    .io_spriteXPosition_25(graphicEngineVGA_io_spriteXPosition_25),
    .io_spriteXPosition_26(graphicEngineVGA_io_spriteXPosition_26),
    .io_spriteXPosition_27(graphicEngineVGA_io_spriteXPosition_27),
    .io_spriteXPosition_28(graphicEngineVGA_io_spriteXPosition_28),
    .io_spriteXPosition_29(graphicEngineVGA_io_spriteXPosition_29),
    .io_spriteXPosition_30(graphicEngineVGA_io_spriteXPosition_30),
    .io_spriteXPosition_31(graphicEngineVGA_io_spriteXPosition_31),
    .io_spriteXPosition_32(graphicEngineVGA_io_spriteXPosition_32),
    .io_spriteXPosition_33(graphicEngineVGA_io_spriteXPosition_33),
    .io_spriteXPosition_34(graphicEngineVGA_io_spriteXPosition_34),
    .io_spriteXPosition_35(graphicEngineVGA_io_spriteXPosition_35),
    .io_spriteXPosition_36(graphicEngineVGA_io_spriteXPosition_36),
    .io_spriteXPosition_37(graphicEngineVGA_io_spriteXPosition_37),
    .io_spriteXPosition_38(graphicEngineVGA_io_spriteXPosition_38),
    .io_spriteXPosition_39(graphicEngineVGA_io_spriteXPosition_39),
    .io_spriteXPosition_40(graphicEngineVGA_io_spriteXPosition_40),
    .io_spriteXPosition_41(graphicEngineVGA_io_spriteXPosition_41),
    .io_spriteXPosition_42(graphicEngineVGA_io_spriteXPosition_42),
    .io_spriteXPosition_43(graphicEngineVGA_io_spriteXPosition_43),
    .io_spriteXPosition_44(graphicEngineVGA_io_spriteXPosition_44),
    .io_spriteXPosition_45(graphicEngineVGA_io_spriteXPosition_45),
    .io_spriteXPosition_46(graphicEngineVGA_io_spriteXPosition_46),
    .io_spriteXPosition_47(graphicEngineVGA_io_spriteXPosition_47),
    .io_spriteXPosition_48(graphicEngineVGA_io_spriteXPosition_48),
    .io_spriteXPosition_49(graphicEngineVGA_io_spriteXPosition_49),
    .io_spriteXPosition_50(graphicEngineVGA_io_spriteXPosition_50),
    .io_spriteXPosition_51(graphicEngineVGA_io_spriteXPosition_51),
    .io_spriteXPosition_52(graphicEngineVGA_io_spriteXPosition_52),
    .io_spriteXPosition_53(graphicEngineVGA_io_spriteXPosition_53),
    .io_spriteXPosition_54(graphicEngineVGA_io_spriteXPosition_54),
    .io_spriteXPosition_55(graphicEngineVGA_io_spriteXPosition_55),
    .io_spriteXPosition_56(graphicEngineVGA_io_spriteXPosition_56),
    .io_spriteXPosition_57(graphicEngineVGA_io_spriteXPosition_57),
    .io_spriteXPosition_58(graphicEngineVGA_io_spriteXPosition_58),
    .io_spriteXPosition_59(graphicEngineVGA_io_spriteXPosition_59),
    .io_spriteXPosition_60(graphicEngineVGA_io_spriteXPosition_60),
    .io_spriteXPosition_61(graphicEngineVGA_io_spriteXPosition_61),
    .io_spriteXPosition_62(graphicEngineVGA_io_spriteXPosition_62),
    .io_spriteXPosition_63(graphicEngineVGA_io_spriteXPosition_63),
    .io_spriteYPosition_3(graphicEngineVGA_io_spriteYPosition_3),
    .io_spriteYPosition_7(graphicEngineVGA_io_spriteYPosition_7),
    .io_spriteYPosition_8(graphicEngineVGA_io_spriteYPosition_8),
    .io_spriteYPosition_9(graphicEngineVGA_io_spriteYPosition_9),
    .io_spriteYPosition_10(graphicEngineVGA_io_spriteYPosition_10),
    .io_spriteYPosition_11(graphicEngineVGA_io_spriteYPosition_11),
    .io_spriteYPosition_12(graphicEngineVGA_io_spriteYPosition_12),
    .io_spriteYPosition_13(graphicEngineVGA_io_spriteYPosition_13),
    .io_spriteYPosition_14(graphicEngineVGA_io_spriteYPosition_14),
    .io_spriteYPosition_16(graphicEngineVGA_io_spriteYPosition_16),
    .io_spriteYPosition_17(graphicEngineVGA_io_spriteYPosition_17),
    .io_spriteYPosition_18(graphicEngineVGA_io_spriteYPosition_18),
    .io_spriteYPosition_19(graphicEngineVGA_io_spriteYPosition_19),
    .io_spriteYPosition_20(graphicEngineVGA_io_spriteYPosition_20),
    .io_spriteYPosition_21(graphicEngineVGA_io_spriteYPosition_21),
    .io_spriteYPosition_22(graphicEngineVGA_io_spriteYPosition_22),
    .io_spriteYPosition_23(graphicEngineVGA_io_spriteYPosition_23),
    .io_spriteYPosition_24(graphicEngineVGA_io_spriteYPosition_24),
    .io_spriteYPosition_25(graphicEngineVGA_io_spriteYPosition_25),
    .io_spriteYPosition_26(graphicEngineVGA_io_spriteYPosition_26),
    .io_spriteYPosition_27(graphicEngineVGA_io_spriteYPosition_27),
    .io_spriteYPosition_28(graphicEngineVGA_io_spriteYPosition_28),
    .io_spriteYPosition_29(graphicEngineVGA_io_spriteYPosition_29),
    .io_spriteYPosition_30(graphicEngineVGA_io_spriteYPosition_30),
    .io_spriteYPosition_31(graphicEngineVGA_io_spriteYPosition_31),
    .io_spriteYPosition_32(graphicEngineVGA_io_spriteYPosition_32),
    .io_spriteYPosition_33(graphicEngineVGA_io_spriteYPosition_33),
    .io_spriteYPosition_34(graphicEngineVGA_io_spriteYPosition_34),
    .io_spriteYPosition_35(graphicEngineVGA_io_spriteYPosition_35),
    .io_spriteYPosition_36(graphicEngineVGA_io_spriteYPosition_36),
    .io_spriteYPosition_37(graphicEngineVGA_io_spriteYPosition_37),
    .io_spriteYPosition_38(graphicEngineVGA_io_spriteYPosition_38),
    .io_spriteYPosition_39(graphicEngineVGA_io_spriteYPosition_39),
    .io_spriteYPosition_40(graphicEngineVGA_io_spriteYPosition_40),
    .io_spriteYPosition_41(graphicEngineVGA_io_spriteYPosition_41),
    .io_spriteYPosition_42(graphicEngineVGA_io_spriteYPosition_42),
    .io_spriteYPosition_43(graphicEngineVGA_io_spriteYPosition_43),
    .io_spriteYPosition_44(graphicEngineVGA_io_spriteYPosition_44),
    .io_spriteYPosition_45(graphicEngineVGA_io_spriteYPosition_45),
    .io_spriteYPosition_46(graphicEngineVGA_io_spriteYPosition_46),
    .io_spriteYPosition_47(graphicEngineVGA_io_spriteYPosition_47),
    .io_spriteYPosition_48(graphicEngineVGA_io_spriteYPosition_48),
    .io_spriteYPosition_49(graphicEngineVGA_io_spriteYPosition_49),
    .io_spriteYPosition_50(graphicEngineVGA_io_spriteYPosition_50),
    .io_spriteYPosition_51(graphicEngineVGA_io_spriteYPosition_51),
    .io_spriteYPosition_52(graphicEngineVGA_io_spriteYPosition_52),
    .io_spriteYPosition_53(graphicEngineVGA_io_spriteYPosition_53),
    .io_spriteYPosition_54(graphicEngineVGA_io_spriteYPosition_54),
    .io_spriteYPosition_55(graphicEngineVGA_io_spriteYPosition_55),
    .io_spriteYPosition_56(graphicEngineVGA_io_spriteYPosition_56),
    .io_spriteYPosition_57(graphicEngineVGA_io_spriteYPosition_57),
    .io_spriteYPosition_58(graphicEngineVGA_io_spriteYPosition_58),
    .io_spriteYPosition_59(graphicEngineVGA_io_spriteYPosition_59),
    .io_spriteYPosition_60(graphicEngineVGA_io_spriteYPosition_60),
    .io_spriteYPosition_61(graphicEngineVGA_io_spriteYPosition_61),
    .io_spriteYPosition_62(graphicEngineVGA_io_spriteYPosition_62),
    .io_spriteYPosition_63(graphicEngineVGA_io_spriteYPosition_63),
    .io_spriteVisible_3(graphicEngineVGA_io_spriteVisible_3),
    .io_spriteVisible_4(graphicEngineVGA_io_spriteVisible_4),
    .io_spriteVisible_5(graphicEngineVGA_io_spriteVisible_5),
    .io_spriteVisible_6(graphicEngineVGA_io_spriteVisible_6),
    .io_spriteVisible_7(graphicEngineVGA_io_spriteVisible_7),
    .io_spriteVisible_8(graphicEngineVGA_io_spriteVisible_8),
    .io_spriteVisible_9(graphicEngineVGA_io_spriteVisible_9),
    .io_spriteVisible_10(graphicEngineVGA_io_spriteVisible_10),
    .io_spriteVisible_11(graphicEngineVGA_io_spriteVisible_11),
    .io_spriteVisible_12(graphicEngineVGA_io_spriteVisible_12),
    .io_spriteVisible_13(graphicEngineVGA_io_spriteVisible_13),
    .io_spriteVisible_14(graphicEngineVGA_io_spriteVisible_14),
    .io_spriteVisible_15(graphicEngineVGA_io_spriteVisible_15),
    .io_spriteVisible_16(graphicEngineVGA_io_spriteVisible_16),
    .io_spriteVisible_17(graphicEngineVGA_io_spriteVisible_17),
    .io_spriteVisible_18(graphicEngineVGA_io_spriteVisible_18),
    .io_spriteVisible_19(graphicEngineVGA_io_spriteVisible_19),
    .io_spriteVisible_20(graphicEngineVGA_io_spriteVisible_20),
    .io_spriteVisible_21(graphicEngineVGA_io_spriteVisible_21),
    .io_spriteVisible_22(graphicEngineVGA_io_spriteVisible_22),
    .io_spriteVisible_23(graphicEngineVGA_io_spriteVisible_23),
    .io_spriteVisible_24(graphicEngineVGA_io_spriteVisible_24),
    .io_spriteVisible_25(graphicEngineVGA_io_spriteVisible_25),
    .io_spriteVisible_26(graphicEngineVGA_io_spriteVisible_26),
    .io_spriteVisible_27(graphicEngineVGA_io_spriteVisible_27),
    .io_spriteVisible_28(graphicEngineVGA_io_spriteVisible_28),
    .io_spriteVisible_29(graphicEngineVGA_io_spriteVisible_29),
    .io_spriteVisible_30(graphicEngineVGA_io_spriteVisible_30),
    .io_spriteVisible_31(graphicEngineVGA_io_spriteVisible_31),
    .io_spriteVisible_32(graphicEngineVGA_io_spriteVisible_32),
    .io_spriteVisible_33(graphicEngineVGA_io_spriteVisible_33),
    .io_spriteVisible_34(graphicEngineVGA_io_spriteVisible_34),
    .io_spriteVisible_35(graphicEngineVGA_io_spriteVisible_35),
    .io_spriteVisible_36(graphicEngineVGA_io_spriteVisible_36),
    .io_spriteVisible_37(graphicEngineVGA_io_spriteVisible_37),
    .io_spriteVisible_38(graphicEngineVGA_io_spriteVisible_38),
    .io_spriteVisible_39(graphicEngineVGA_io_spriteVisible_39),
    .io_spriteVisible_40(graphicEngineVGA_io_spriteVisible_40),
    .io_spriteVisible_41(graphicEngineVGA_io_spriteVisible_41),
    .io_spriteVisible_42(graphicEngineVGA_io_spriteVisible_42),
    .io_spriteVisible_43(graphicEngineVGA_io_spriteVisible_43),
    .io_spriteVisible_44(graphicEngineVGA_io_spriteVisible_44),
    .io_spriteVisible_45(graphicEngineVGA_io_spriteVisible_45),
    .io_spriteVisible_46(graphicEngineVGA_io_spriteVisible_46),
    .io_spriteVisible_47(graphicEngineVGA_io_spriteVisible_47),
    .io_spriteVisible_48(graphicEngineVGA_io_spriteVisible_48),
    .io_spriteVisible_49(graphicEngineVGA_io_spriteVisible_49),
    .io_spriteVisible_50(graphicEngineVGA_io_spriteVisible_50),
    .io_spriteVisible_51(graphicEngineVGA_io_spriteVisible_51),
    .io_spriteVisible_52(graphicEngineVGA_io_spriteVisible_52),
    .io_spriteVisible_53(graphicEngineVGA_io_spriteVisible_53),
    .io_spriteVisible_54(graphicEngineVGA_io_spriteVisible_54),
    .io_spriteVisible_55(graphicEngineVGA_io_spriteVisible_55),
    .io_spriteVisible_56(graphicEngineVGA_io_spriteVisible_56),
    .io_spriteVisible_57(graphicEngineVGA_io_spriteVisible_57),
    .io_spriteVisible_58(graphicEngineVGA_io_spriteVisible_58),
    .io_spriteVisible_59(graphicEngineVGA_io_spriteVisible_59),
    .io_spriteVisible_60(graphicEngineVGA_io_spriteVisible_60),
    .io_spriteVisible_61(graphicEngineVGA_io_spriteVisible_61),
    .io_spriteVisible_62(graphicEngineVGA_io_spriteVisible_62),
    .io_spriteVisible_63(graphicEngineVGA_io_spriteVisible_63),
    .io_spriteScaleUpHorizontal_16(graphicEngineVGA_io_spriteScaleUpHorizontal_16),
    .io_spriteScaleUpHorizontal_17(graphicEngineVGA_io_spriteScaleUpHorizontal_17),
    .io_spriteScaleUpHorizontal_18(graphicEngineVGA_io_spriteScaleUpHorizontal_18),
    .io_spriteScaleUpHorizontal_19(graphicEngineVGA_io_spriteScaleUpHorizontal_19),
    .io_spriteScaleUpHorizontal_20(graphicEngineVGA_io_spriteScaleUpHorizontal_20),
    .io_spriteScaleUpHorizontal_21(graphicEngineVGA_io_spriteScaleUpHorizontal_21),
    .io_spriteScaleUpHorizontal_22(graphicEngineVGA_io_spriteScaleUpHorizontal_22),
    .io_spriteScaleUpHorizontal_23(graphicEngineVGA_io_spriteScaleUpHorizontal_23),
    .io_spriteScaleUpHorizontal_24(graphicEngineVGA_io_spriteScaleUpHorizontal_24),
    .io_spriteScaleUpHorizontal_25(graphicEngineVGA_io_spriteScaleUpHorizontal_25),
    .io_spriteScaleUpHorizontal_26(graphicEngineVGA_io_spriteScaleUpHorizontal_26),
    .io_spriteScaleUpHorizontal_27(graphicEngineVGA_io_spriteScaleUpHorizontal_27),
    .io_spriteScaleUpHorizontal_28(graphicEngineVGA_io_spriteScaleUpHorizontal_28),
    .io_spriteScaleUpHorizontal_29(graphicEngineVGA_io_spriteScaleUpHorizontal_29),
    .io_spriteScaleUpHorizontal_30(graphicEngineVGA_io_spriteScaleUpHorizontal_30),
    .io_spriteScaleUpHorizontal_31(graphicEngineVGA_io_spriteScaleUpHorizontal_31),
    .io_spriteScaleUpHorizontal_32(graphicEngineVGA_io_spriteScaleUpHorizontal_32),
    .io_spriteScaleUpHorizontal_33(graphicEngineVGA_io_spriteScaleUpHorizontal_33),
    .io_spriteScaleUpHorizontal_34(graphicEngineVGA_io_spriteScaleUpHorizontal_34),
    .io_spriteScaleUpHorizontal_35(graphicEngineVGA_io_spriteScaleUpHorizontal_35),
    .io_spriteScaleUpHorizontal_36(graphicEngineVGA_io_spriteScaleUpHorizontal_36),
    .io_spriteScaleUpHorizontal_37(graphicEngineVGA_io_spriteScaleUpHorizontal_37),
    .io_spriteScaleUpHorizontal_38(graphicEngineVGA_io_spriteScaleUpHorizontal_38),
    .io_spriteScaleUpHorizontal_39(graphicEngineVGA_io_spriteScaleUpHorizontal_39),
    .io_spriteScaleUpHorizontal_40(graphicEngineVGA_io_spriteScaleUpHorizontal_40),
    .io_spriteScaleUpHorizontal_41(graphicEngineVGA_io_spriteScaleUpHorizontal_41),
    .io_spriteScaleUpHorizontal_42(graphicEngineVGA_io_spriteScaleUpHorizontal_42),
    .io_spriteScaleUpHorizontal_43(graphicEngineVGA_io_spriteScaleUpHorizontal_43),
    .io_spriteScaleUpHorizontal_44(graphicEngineVGA_io_spriteScaleUpHorizontal_44),
    .io_spriteScaleUpHorizontal_45(graphicEngineVGA_io_spriteScaleUpHorizontal_45),
    .io_spriteScaleUpHorizontal_58(graphicEngineVGA_io_spriteScaleUpHorizontal_58),
    .io_spriteScaleUpHorizontal_59(graphicEngineVGA_io_spriteScaleUpHorizontal_59),
    .io_spriteScaleUpHorizontal_60(graphicEngineVGA_io_spriteScaleUpHorizontal_60),
    .io_spriteScaleUpVertical_16(graphicEngineVGA_io_spriteScaleUpVertical_16),
    .io_spriteScaleUpVertical_17(graphicEngineVGA_io_spriteScaleUpVertical_17),
    .io_spriteScaleUpVertical_18(graphicEngineVGA_io_spriteScaleUpVertical_18),
    .io_spriteScaleUpVertical_19(graphicEngineVGA_io_spriteScaleUpVertical_19),
    .io_spriteScaleUpVertical_20(graphicEngineVGA_io_spriteScaleUpVertical_20),
    .io_spriteScaleUpVertical_21(graphicEngineVGA_io_spriteScaleUpVertical_21),
    .io_spriteScaleUpVertical_22(graphicEngineVGA_io_spriteScaleUpVertical_22),
    .io_spriteScaleUpVertical_23(graphicEngineVGA_io_spriteScaleUpVertical_23),
    .io_spriteScaleUpVertical_24(graphicEngineVGA_io_spriteScaleUpVertical_24),
    .io_spriteScaleUpVertical_25(graphicEngineVGA_io_spriteScaleUpVertical_25),
    .io_spriteScaleUpVertical_26(graphicEngineVGA_io_spriteScaleUpVertical_26),
    .io_spriteScaleUpVertical_27(graphicEngineVGA_io_spriteScaleUpVertical_27),
    .io_spriteScaleUpVertical_28(graphicEngineVGA_io_spriteScaleUpVertical_28),
    .io_spriteScaleUpVertical_29(graphicEngineVGA_io_spriteScaleUpVertical_29),
    .io_spriteScaleUpVertical_30(graphicEngineVGA_io_spriteScaleUpVertical_30),
    .io_spriteScaleUpVertical_31(graphicEngineVGA_io_spriteScaleUpVertical_31),
    .io_spriteScaleUpVertical_32(graphicEngineVGA_io_spriteScaleUpVertical_32),
    .io_spriteScaleUpVertical_33(graphicEngineVGA_io_spriteScaleUpVertical_33),
    .io_spriteScaleUpVertical_34(graphicEngineVGA_io_spriteScaleUpVertical_34),
    .io_spriteScaleUpVertical_35(graphicEngineVGA_io_spriteScaleUpVertical_35),
    .io_spriteScaleUpVertical_36(graphicEngineVGA_io_spriteScaleUpVertical_36),
    .io_spriteScaleUpVertical_37(graphicEngineVGA_io_spriteScaleUpVertical_37),
    .io_spriteScaleUpVertical_38(graphicEngineVGA_io_spriteScaleUpVertical_38),
    .io_spriteScaleUpVertical_39(graphicEngineVGA_io_spriteScaleUpVertical_39),
    .io_spriteScaleUpVertical_40(graphicEngineVGA_io_spriteScaleUpVertical_40),
    .io_spriteScaleUpVertical_41(graphicEngineVGA_io_spriteScaleUpVertical_41),
    .io_spriteScaleUpVertical_42(graphicEngineVGA_io_spriteScaleUpVertical_42),
    .io_spriteScaleUpVertical_43(graphicEngineVGA_io_spriteScaleUpVertical_43),
    .io_spriteScaleUpVertical_44(graphicEngineVGA_io_spriteScaleUpVertical_44),
    .io_spriteScaleUpVertical_45(graphicEngineVGA_io_spriteScaleUpVertical_45),
    .io_spriteScaleUpVertical_58(graphicEngineVGA_io_spriteScaleUpVertical_58),
    .io_spriteScaleUpVertical_59(graphicEngineVGA_io_spriteScaleUpVertical_59),
    .io_spriteScaleUpVertical_60(graphicEngineVGA_io_spriteScaleUpVertical_60),
    .io_viewBoxX(graphicEngineVGA_io_viewBoxX),
    .io_viewBoxY(graphicEngineVGA_io_viewBoxY),
    .io_newFrame(graphicEngineVGA_io_newFrame),
    .io_frameUpdateDone(graphicEngineVGA_io_frameUpdateDone),
    .io_missingFrameError(graphicEngineVGA_io_missingFrameError),
    .io_viewBoxOutOfRangeError(graphicEngineVGA_io_viewBoxOutOfRangeError),
    .io_vgaRed(graphicEngineVGA_io_vgaRed),
    .io_vgaBlue(graphicEngineVGA_io_vgaBlue),
    .io_vgaGreen(graphicEngineVGA_io_vgaGreen),
    .io_Hsync(graphicEngineVGA_io_Hsync),
    .io_Vsync(graphicEngineVGA_io_Vsync)
  );
  SoundEngine soundEngine ( // @[\\src\\main\\scala\\GameTop.scala 49:27]
    .clock(soundEngine_clock),
    .reset(soundEngine_reset)
  );
  GameLogic gameLogic ( // @[\\src\\main\\scala\\GameTop.scala 53:25]
    .clock(gameLogic_clock),
    .reset(gameLogic_reset),
    .io_btnC(gameLogic_io_btnC),
    .io_btnU(gameLogic_io_btnU),
    .io_btnL(gameLogic_io_btnL),
    .io_btnR(gameLogic_io_btnR),
    .io_btnD(gameLogic_io_btnD),
    .io_spriteXPosition_3(gameLogic_io_spriteXPosition_3),
    .io_spriteXPosition_7(gameLogic_io_spriteXPosition_7),
    .io_spriteXPosition_8(gameLogic_io_spriteXPosition_8),
    .io_spriteXPosition_9(gameLogic_io_spriteXPosition_9),
    .io_spriteXPosition_10(gameLogic_io_spriteXPosition_10),
    .io_spriteXPosition_11(gameLogic_io_spriteXPosition_11),
    .io_spriteXPosition_12(gameLogic_io_spriteXPosition_12),
    .io_spriteXPosition_13(gameLogic_io_spriteXPosition_13),
    .io_spriteXPosition_14(gameLogic_io_spriteXPosition_14),
    .io_spriteXPosition_16(gameLogic_io_spriteXPosition_16),
    .io_spriteXPosition_17(gameLogic_io_spriteXPosition_17),
    .io_spriteXPosition_18(gameLogic_io_spriteXPosition_18),
    .io_spriteXPosition_19(gameLogic_io_spriteXPosition_19),
    .io_spriteXPosition_20(gameLogic_io_spriteXPosition_20),
    .io_spriteXPosition_21(gameLogic_io_spriteXPosition_21),
    .io_spriteXPosition_22(gameLogic_io_spriteXPosition_22),
    .io_spriteXPosition_23(gameLogic_io_spriteXPosition_23),
    .io_spriteXPosition_24(gameLogic_io_spriteXPosition_24),
    .io_spriteXPosition_25(gameLogic_io_spriteXPosition_25),
    .io_spriteXPosition_26(gameLogic_io_spriteXPosition_26),
    .io_spriteXPosition_27(gameLogic_io_spriteXPosition_27),
    .io_spriteXPosition_28(gameLogic_io_spriteXPosition_28),
    .io_spriteXPosition_29(gameLogic_io_spriteXPosition_29),
    .io_spriteXPosition_30(gameLogic_io_spriteXPosition_30),
    .io_spriteXPosition_31(gameLogic_io_spriteXPosition_31),
    .io_spriteXPosition_32(gameLogic_io_spriteXPosition_32),
    .io_spriteXPosition_33(gameLogic_io_spriteXPosition_33),
    .io_spriteXPosition_34(gameLogic_io_spriteXPosition_34),
    .io_spriteXPosition_35(gameLogic_io_spriteXPosition_35),
    .io_spriteXPosition_36(gameLogic_io_spriteXPosition_36),
    .io_spriteXPosition_37(gameLogic_io_spriteXPosition_37),
    .io_spriteXPosition_38(gameLogic_io_spriteXPosition_38),
    .io_spriteXPosition_39(gameLogic_io_spriteXPosition_39),
    .io_spriteXPosition_40(gameLogic_io_spriteXPosition_40),
    .io_spriteXPosition_41(gameLogic_io_spriteXPosition_41),
    .io_spriteXPosition_42(gameLogic_io_spriteXPosition_42),
    .io_spriteXPosition_43(gameLogic_io_spriteXPosition_43),
    .io_spriteXPosition_44(gameLogic_io_spriteXPosition_44),
    .io_spriteXPosition_45(gameLogic_io_spriteXPosition_45),
    .io_spriteXPosition_46(gameLogic_io_spriteXPosition_46),
    .io_spriteXPosition_47(gameLogic_io_spriteXPosition_47),
    .io_spriteXPosition_48(gameLogic_io_spriteXPosition_48),
    .io_spriteXPosition_49(gameLogic_io_spriteXPosition_49),
    .io_spriteXPosition_50(gameLogic_io_spriteXPosition_50),
    .io_spriteXPosition_51(gameLogic_io_spriteXPosition_51),
    .io_spriteXPosition_52(gameLogic_io_spriteXPosition_52),
    .io_spriteXPosition_53(gameLogic_io_spriteXPosition_53),
    .io_spriteXPosition_54(gameLogic_io_spriteXPosition_54),
    .io_spriteXPosition_55(gameLogic_io_spriteXPosition_55),
    .io_spriteXPosition_56(gameLogic_io_spriteXPosition_56),
    .io_spriteXPosition_57(gameLogic_io_spriteXPosition_57),
    .io_spriteXPosition_58(gameLogic_io_spriteXPosition_58),
    .io_spriteXPosition_59(gameLogic_io_spriteXPosition_59),
    .io_spriteXPosition_60(gameLogic_io_spriteXPosition_60),
    .io_spriteXPosition_61(gameLogic_io_spriteXPosition_61),
    .io_spriteXPosition_62(gameLogic_io_spriteXPosition_62),
    .io_spriteXPosition_63(gameLogic_io_spriteXPosition_63),
    .io_spriteYPosition_3(gameLogic_io_spriteYPosition_3),
    .io_spriteYPosition_7(gameLogic_io_spriteYPosition_7),
    .io_spriteYPosition_8(gameLogic_io_spriteYPosition_8),
    .io_spriteYPosition_9(gameLogic_io_spriteYPosition_9),
    .io_spriteYPosition_10(gameLogic_io_spriteYPosition_10),
    .io_spriteYPosition_11(gameLogic_io_spriteYPosition_11),
    .io_spriteYPosition_12(gameLogic_io_spriteYPosition_12),
    .io_spriteYPosition_13(gameLogic_io_spriteYPosition_13),
    .io_spriteYPosition_14(gameLogic_io_spriteYPosition_14),
    .io_spriteYPosition_16(gameLogic_io_spriteYPosition_16),
    .io_spriteYPosition_17(gameLogic_io_spriteYPosition_17),
    .io_spriteYPosition_18(gameLogic_io_spriteYPosition_18),
    .io_spriteYPosition_19(gameLogic_io_spriteYPosition_19),
    .io_spriteYPosition_20(gameLogic_io_spriteYPosition_20),
    .io_spriteYPosition_21(gameLogic_io_spriteYPosition_21),
    .io_spriteYPosition_22(gameLogic_io_spriteYPosition_22),
    .io_spriteYPosition_23(gameLogic_io_spriteYPosition_23),
    .io_spriteYPosition_24(gameLogic_io_spriteYPosition_24),
    .io_spriteYPosition_25(gameLogic_io_spriteYPosition_25),
    .io_spriteYPosition_26(gameLogic_io_spriteYPosition_26),
    .io_spriteYPosition_27(gameLogic_io_spriteYPosition_27),
    .io_spriteYPosition_28(gameLogic_io_spriteYPosition_28),
    .io_spriteYPosition_29(gameLogic_io_spriteYPosition_29),
    .io_spriteYPosition_30(gameLogic_io_spriteYPosition_30),
    .io_spriteYPosition_31(gameLogic_io_spriteYPosition_31),
    .io_spriteYPosition_32(gameLogic_io_spriteYPosition_32),
    .io_spriteYPosition_33(gameLogic_io_spriteYPosition_33),
    .io_spriteYPosition_34(gameLogic_io_spriteYPosition_34),
    .io_spriteYPosition_35(gameLogic_io_spriteYPosition_35),
    .io_spriteYPosition_36(gameLogic_io_spriteYPosition_36),
    .io_spriteYPosition_37(gameLogic_io_spriteYPosition_37),
    .io_spriteYPosition_38(gameLogic_io_spriteYPosition_38),
    .io_spriteYPosition_39(gameLogic_io_spriteYPosition_39),
    .io_spriteYPosition_40(gameLogic_io_spriteYPosition_40),
    .io_spriteYPosition_41(gameLogic_io_spriteYPosition_41),
    .io_spriteYPosition_42(gameLogic_io_spriteYPosition_42),
    .io_spriteYPosition_43(gameLogic_io_spriteYPosition_43),
    .io_spriteYPosition_44(gameLogic_io_spriteYPosition_44),
    .io_spriteYPosition_45(gameLogic_io_spriteYPosition_45),
    .io_spriteYPosition_46(gameLogic_io_spriteYPosition_46),
    .io_spriteYPosition_47(gameLogic_io_spriteYPosition_47),
    .io_spriteYPosition_48(gameLogic_io_spriteYPosition_48),
    .io_spriteYPosition_49(gameLogic_io_spriteYPosition_49),
    .io_spriteYPosition_50(gameLogic_io_spriteYPosition_50),
    .io_spriteYPosition_51(gameLogic_io_spriteYPosition_51),
    .io_spriteYPosition_52(gameLogic_io_spriteYPosition_52),
    .io_spriteYPosition_53(gameLogic_io_spriteYPosition_53),
    .io_spriteYPosition_54(gameLogic_io_spriteYPosition_54),
    .io_spriteYPosition_55(gameLogic_io_spriteYPosition_55),
    .io_spriteYPosition_56(gameLogic_io_spriteYPosition_56),
    .io_spriteYPosition_57(gameLogic_io_spriteYPosition_57),
    .io_spriteYPosition_58(gameLogic_io_spriteYPosition_58),
    .io_spriteYPosition_59(gameLogic_io_spriteYPosition_59),
    .io_spriteYPosition_60(gameLogic_io_spriteYPosition_60),
    .io_spriteYPosition_61(gameLogic_io_spriteYPosition_61),
    .io_spriteYPosition_62(gameLogic_io_spriteYPosition_62),
    .io_spriteYPosition_63(gameLogic_io_spriteYPosition_63),
    .io_spriteVisible_3(gameLogic_io_spriteVisible_3),
    .io_spriteVisible_4(gameLogic_io_spriteVisible_4),
    .io_spriteVisible_5(gameLogic_io_spriteVisible_5),
    .io_spriteVisible_6(gameLogic_io_spriteVisible_6),
    .io_spriteVisible_7(gameLogic_io_spriteVisible_7),
    .io_spriteVisible_8(gameLogic_io_spriteVisible_8),
    .io_spriteVisible_9(gameLogic_io_spriteVisible_9),
    .io_spriteVisible_10(gameLogic_io_spriteVisible_10),
    .io_spriteVisible_11(gameLogic_io_spriteVisible_11),
    .io_spriteVisible_12(gameLogic_io_spriteVisible_12),
    .io_spriteVisible_13(gameLogic_io_spriteVisible_13),
    .io_spriteVisible_14(gameLogic_io_spriteVisible_14),
    .io_spriteVisible_15(gameLogic_io_spriteVisible_15),
    .io_spriteVisible_16(gameLogic_io_spriteVisible_16),
    .io_spriteVisible_17(gameLogic_io_spriteVisible_17),
    .io_spriteVisible_18(gameLogic_io_spriteVisible_18),
    .io_spriteVisible_19(gameLogic_io_spriteVisible_19),
    .io_spriteVisible_20(gameLogic_io_spriteVisible_20),
    .io_spriteVisible_21(gameLogic_io_spriteVisible_21),
    .io_spriteVisible_22(gameLogic_io_spriteVisible_22),
    .io_spriteVisible_23(gameLogic_io_spriteVisible_23),
    .io_spriteVisible_24(gameLogic_io_spriteVisible_24),
    .io_spriteVisible_25(gameLogic_io_spriteVisible_25),
    .io_spriteVisible_26(gameLogic_io_spriteVisible_26),
    .io_spriteVisible_27(gameLogic_io_spriteVisible_27),
    .io_spriteVisible_28(gameLogic_io_spriteVisible_28),
    .io_spriteVisible_29(gameLogic_io_spriteVisible_29),
    .io_spriteVisible_30(gameLogic_io_spriteVisible_30),
    .io_spriteVisible_31(gameLogic_io_spriteVisible_31),
    .io_spriteVisible_32(gameLogic_io_spriteVisible_32),
    .io_spriteVisible_33(gameLogic_io_spriteVisible_33),
    .io_spriteVisible_34(gameLogic_io_spriteVisible_34),
    .io_spriteVisible_35(gameLogic_io_spriteVisible_35),
    .io_spriteVisible_36(gameLogic_io_spriteVisible_36),
    .io_spriteVisible_37(gameLogic_io_spriteVisible_37),
    .io_spriteVisible_38(gameLogic_io_spriteVisible_38),
    .io_spriteVisible_39(gameLogic_io_spriteVisible_39),
    .io_spriteVisible_40(gameLogic_io_spriteVisible_40),
    .io_spriteVisible_41(gameLogic_io_spriteVisible_41),
    .io_spriteVisible_42(gameLogic_io_spriteVisible_42),
    .io_spriteVisible_43(gameLogic_io_spriteVisible_43),
    .io_spriteVisible_44(gameLogic_io_spriteVisible_44),
    .io_spriteVisible_45(gameLogic_io_spriteVisible_45),
    .io_spriteVisible_46(gameLogic_io_spriteVisible_46),
    .io_spriteVisible_47(gameLogic_io_spriteVisible_47),
    .io_spriteVisible_48(gameLogic_io_spriteVisible_48),
    .io_spriteVisible_49(gameLogic_io_spriteVisible_49),
    .io_spriteVisible_50(gameLogic_io_spriteVisible_50),
    .io_spriteVisible_51(gameLogic_io_spriteVisible_51),
    .io_spriteVisible_52(gameLogic_io_spriteVisible_52),
    .io_spriteVisible_53(gameLogic_io_spriteVisible_53),
    .io_spriteVisible_54(gameLogic_io_spriteVisible_54),
    .io_spriteVisible_55(gameLogic_io_spriteVisible_55),
    .io_spriteVisible_56(gameLogic_io_spriteVisible_56),
    .io_spriteVisible_57(gameLogic_io_spriteVisible_57),
    .io_spriteVisible_58(gameLogic_io_spriteVisible_58),
    .io_spriteVisible_59(gameLogic_io_spriteVisible_59),
    .io_spriteVisible_60(gameLogic_io_spriteVisible_60),
    .io_spriteVisible_61(gameLogic_io_spriteVisible_61),
    .io_spriteVisible_62(gameLogic_io_spriteVisible_62),
    .io_spriteVisible_63(gameLogic_io_spriteVisible_63),
    .io_spriteScaleUpHorizontal_16(gameLogic_io_spriteScaleUpHorizontal_16),
    .io_spriteScaleUpHorizontal_17(gameLogic_io_spriteScaleUpHorizontal_17),
    .io_spriteScaleUpHorizontal_18(gameLogic_io_spriteScaleUpHorizontal_18),
    .io_spriteScaleUpHorizontal_19(gameLogic_io_spriteScaleUpHorizontal_19),
    .io_spriteScaleUpHorizontal_20(gameLogic_io_spriteScaleUpHorizontal_20),
    .io_spriteScaleUpHorizontal_21(gameLogic_io_spriteScaleUpHorizontal_21),
    .io_spriteScaleUpHorizontal_22(gameLogic_io_spriteScaleUpHorizontal_22),
    .io_spriteScaleUpHorizontal_23(gameLogic_io_spriteScaleUpHorizontal_23),
    .io_spriteScaleUpHorizontal_24(gameLogic_io_spriteScaleUpHorizontal_24),
    .io_spriteScaleUpHorizontal_25(gameLogic_io_spriteScaleUpHorizontal_25),
    .io_spriteScaleUpHorizontal_26(gameLogic_io_spriteScaleUpHorizontal_26),
    .io_spriteScaleUpHorizontal_27(gameLogic_io_spriteScaleUpHorizontal_27),
    .io_spriteScaleUpHorizontal_28(gameLogic_io_spriteScaleUpHorizontal_28),
    .io_spriteScaleUpHorizontal_29(gameLogic_io_spriteScaleUpHorizontal_29),
    .io_spriteScaleUpHorizontal_30(gameLogic_io_spriteScaleUpHorizontal_30),
    .io_spriteScaleUpHorizontal_31(gameLogic_io_spriteScaleUpHorizontal_31),
    .io_spriteScaleUpHorizontal_32(gameLogic_io_spriteScaleUpHorizontal_32),
    .io_spriteScaleUpHorizontal_33(gameLogic_io_spriteScaleUpHorizontal_33),
    .io_spriteScaleUpHorizontal_34(gameLogic_io_spriteScaleUpHorizontal_34),
    .io_spriteScaleUpHorizontal_35(gameLogic_io_spriteScaleUpHorizontal_35),
    .io_spriteScaleUpHorizontal_36(gameLogic_io_spriteScaleUpHorizontal_36),
    .io_spriteScaleUpHorizontal_37(gameLogic_io_spriteScaleUpHorizontal_37),
    .io_spriteScaleUpHorizontal_38(gameLogic_io_spriteScaleUpHorizontal_38),
    .io_spriteScaleUpHorizontal_39(gameLogic_io_spriteScaleUpHorizontal_39),
    .io_spriteScaleUpHorizontal_40(gameLogic_io_spriteScaleUpHorizontal_40),
    .io_spriteScaleUpHorizontal_41(gameLogic_io_spriteScaleUpHorizontal_41),
    .io_spriteScaleUpHorizontal_42(gameLogic_io_spriteScaleUpHorizontal_42),
    .io_spriteScaleUpHorizontal_43(gameLogic_io_spriteScaleUpHorizontal_43),
    .io_spriteScaleUpHorizontal_44(gameLogic_io_spriteScaleUpHorizontal_44),
    .io_spriteScaleUpHorizontal_45(gameLogic_io_spriteScaleUpHorizontal_45),
    .io_spriteScaleUpHorizontal_58(gameLogic_io_spriteScaleUpHorizontal_58),
    .io_spriteScaleUpHorizontal_59(gameLogic_io_spriteScaleUpHorizontal_59),
    .io_spriteScaleUpHorizontal_60(gameLogic_io_spriteScaleUpHorizontal_60),
    .io_spriteScaleUpVertical_16(gameLogic_io_spriteScaleUpVertical_16),
    .io_spriteScaleUpVertical_17(gameLogic_io_spriteScaleUpVertical_17),
    .io_spriteScaleUpVertical_18(gameLogic_io_spriteScaleUpVertical_18),
    .io_spriteScaleUpVertical_19(gameLogic_io_spriteScaleUpVertical_19),
    .io_spriteScaleUpVertical_20(gameLogic_io_spriteScaleUpVertical_20),
    .io_spriteScaleUpVertical_21(gameLogic_io_spriteScaleUpVertical_21),
    .io_spriteScaleUpVertical_22(gameLogic_io_spriteScaleUpVertical_22),
    .io_spriteScaleUpVertical_23(gameLogic_io_spriteScaleUpVertical_23),
    .io_spriteScaleUpVertical_24(gameLogic_io_spriteScaleUpVertical_24),
    .io_spriteScaleUpVertical_25(gameLogic_io_spriteScaleUpVertical_25),
    .io_spriteScaleUpVertical_26(gameLogic_io_spriteScaleUpVertical_26),
    .io_spriteScaleUpVertical_27(gameLogic_io_spriteScaleUpVertical_27),
    .io_spriteScaleUpVertical_28(gameLogic_io_spriteScaleUpVertical_28),
    .io_spriteScaleUpVertical_29(gameLogic_io_spriteScaleUpVertical_29),
    .io_spriteScaleUpVertical_30(gameLogic_io_spriteScaleUpVertical_30),
    .io_spriteScaleUpVertical_31(gameLogic_io_spriteScaleUpVertical_31),
    .io_spriteScaleUpVertical_32(gameLogic_io_spriteScaleUpVertical_32),
    .io_spriteScaleUpVertical_33(gameLogic_io_spriteScaleUpVertical_33),
    .io_spriteScaleUpVertical_34(gameLogic_io_spriteScaleUpVertical_34),
    .io_spriteScaleUpVertical_35(gameLogic_io_spriteScaleUpVertical_35),
    .io_spriteScaleUpVertical_36(gameLogic_io_spriteScaleUpVertical_36),
    .io_spriteScaleUpVertical_37(gameLogic_io_spriteScaleUpVertical_37),
    .io_spriteScaleUpVertical_38(gameLogic_io_spriteScaleUpVertical_38),
    .io_spriteScaleUpVertical_39(gameLogic_io_spriteScaleUpVertical_39),
    .io_spriteScaleUpVertical_40(gameLogic_io_spriteScaleUpVertical_40),
    .io_spriteScaleUpVertical_41(gameLogic_io_spriteScaleUpVertical_41),
    .io_spriteScaleUpVertical_42(gameLogic_io_spriteScaleUpVertical_42),
    .io_spriteScaleUpVertical_43(gameLogic_io_spriteScaleUpVertical_43),
    .io_spriteScaleUpVertical_44(gameLogic_io_spriteScaleUpVertical_44),
    .io_spriteScaleUpVertical_45(gameLogic_io_spriteScaleUpVertical_45),
    .io_spriteScaleUpVertical_58(gameLogic_io_spriteScaleUpVertical_58),
    .io_spriteScaleUpVertical_59(gameLogic_io_spriteScaleUpVertical_59),
    .io_spriteScaleUpVertical_60(gameLogic_io_spriteScaleUpVertical_60),
    .io_viewBoxX(gameLogic_io_viewBoxX),
    .io_viewBoxY(gameLogic_io_viewBoxY),
    .io_newFrame(gameLogic_io_newFrame),
    .io_frameUpdateDone(gameLogic_io_frameUpdateDone)
  );
  assign io_vgaRed = graphicEngineVGA_io_vgaRed; // @[\\src\\main\\scala\\GameTop.scala 105:13]
  assign io_vgaBlue = graphicEngineVGA_io_vgaBlue; // @[\\src\\main\\scala\\GameTop.scala 107:14]
  assign io_vgaGreen = graphicEngineVGA_io_vgaGreen; // @[\\src\\main\\scala\\GameTop.scala 106:15]
  assign io_Hsync = graphicEngineVGA_io_Hsync; // @[\\src\\main\\scala\\GameTop.scala 108:12]
  assign io_Vsync = graphicEngineVGA_io_Vsync; // @[\\src\\main\\scala\\GameTop.scala 109:12]
  assign io_missingFrameError = graphicEngineVGA_io_missingFrameError; // @[\\src\\main\\scala\\GameTop.scala 120:24]
  assign io_viewBoxOutOfRangeError = graphicEngineVGA_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\GameTop.scala 122:29]
  assign graphicEngineVGA_clock = clock;
  assign graphicEngineVGA_reset = resetReleaseCounter == 22'h3d08ff ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameTop.scala 83:67 84:18 86:18]
  assign graphicEngineVGA_io_spriteXPosition_3 = gameLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_7 = gameLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_8 = gameLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_9 = gameLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_10 = gameLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_11 = gameLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_12 = gameLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_13 = gameLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_14 = gameLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_16 = gameLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_17 = gameLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_18 = gameLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_19 = gameLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_20 = gameLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_21 = gameLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_22 = gameLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_23 = gameLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_24 = gameLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_25 = gameLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_26 = gameLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_27 = gameLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_28 = gameLogic_io_spriteXPosition_28; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_29 = gameLogic_io_spriteXPosition_29; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_30 = gameLogic_io_spriteXPosition_30; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_31 = gameLogic_io_spriteXPosition_31; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_32 = gameLogic_io_spriteXPosition_32; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_33 = gameLogic_io_spriteXPosition_33; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_34 = gameLogic_io_spriteXPosition_34; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_35 = gameLogic_io_spriteXPosition_35; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_36 = gameLogic_io_spriteXPosition_36; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_37 = gameLogic_io_spriteXPosition_37; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_38 = gameLogic_io_spriteXPosition_38; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_39 = gameLogic_io_spriteXPosition_39; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_40 = gameLogic_io_spriteXPosition_40; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_41 = gameLogic_io_spriteXPosition_41; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_42 = gameLogic_io_spriteXPosition_42; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_43 = gameLogic_io_spriteXPosition_43; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_44 = gameLogic_io_spriteXPosition_44; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_45 = gameLogic_io_spriteXPosition_45; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_46 = gameLogic_io_spriteXPosition_46; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_47 = gameLogic_io_spriteXPosition_47; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_48 = gameLogic_io_spriteXPosition_48; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_49 = gameLogic_io_spriteXPosition_49; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_50 = gameLogic_io_spriteXPosition_50; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_51 = gameLogic_io_spriteXPosition_51; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_52 = gameLogic_io_spriteXPosition_52; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_53 = gameLogic_io_spriteXPosition_53; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_54 = gameLogic_io_spriteXPosition_54; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_55 = gameLogic_io_spriteXPosition_55; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_56 = gameLogic_io_spriteXPosition_56; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_57 = gameLogic_io_spriteXPosition_57; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_58 = gameLogic_io_spriteXPosition_58; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_59 = gameLogic_io_spriteXPosition_59; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_60 = gameLogic_io_spriteXPosition_60; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_61 = gameLogic_io_spriteXPosition_61; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_62 = gameLogic_io_spriteXPosition_62; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteXPosition_63 = gameLogic_io_spriteXPosition_63; // @[\\src\\main\\scala\\GameTop.scala 125:39]
  assign graphicEngineVGA_io_spriteYPosition_3 = gameLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_7 = gameLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_8 = gameLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_9 = gameLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_10 = gameLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_11 = gameLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_12 = gameLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_13 = gameLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_14 = gameLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_16 = gameLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_17 = gameLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_18 = gameLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_19 = gameLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_20 = gameLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_21 = gameLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_22 = gameLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_23 = gameLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_24 = gameLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_25 = gameLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_26 = gameLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_27 = gameLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_28 = gameLogic_io_spriteYPosition_28; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_29 = gameLogic_io_spriteYPosition_29; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_30 = gameLogic_io_spriteYPosition_30; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_31 = gameLogic_io_spriteYPosition_31; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_32 = gameLogic_io_spriteYPosition_32; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_33 = gameLogic_io_spriteYPosition_33; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_34 = gameLogic_io_spriteYPosition_34; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_35 = gameLogic_io_spriteYPosition_35; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_36 = gameLogic_io_spriteYPosition_36; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_37 = gameLogic_io_spriteYPosition_37; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_38 = gameLogic_io_spriteYPosition_38; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_39 = gameLogic_io_spriteYPosition_39; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_40 = gameLogic_io_spriteYPosition_40; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_41 = gameLogic_io_spriteYPosition_41; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_42 = gameLogic_io_spriteYPosition_42; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_43 = gameLogic_io_spriteYPosition_43; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_44 = gameLogic_io_spriteYPosition_44; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_45 = gameLogic_io_spriteYPosition_45; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_46 = gameLogic_io_spriteYPosition_46; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_47 = gameLogic_io_spriteYPosition_47; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_48 = gameLogic_io_spriteYPosition_48; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_49 = gameLogic_io_spriteYPosition_49; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_50 = gameLogic_io_spriteYPosition_50; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_51 = gameLogic_io_spriteYPosition_51; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_52 = gameLogic_io_spriteYPosition_52; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_53 = gameLogic_io_spriteYPosition_53; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_54 = gameLogic_io_spriteYPosition_54; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_55 = gameLogic_io_spriteYPosition_55; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_56 = gameLogic_io_spriteYPosition_56; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_57 = gameLogic_io_spriteYPosition_57; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_58 = gameLogic_io_spriteYPosition_58; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_59 = gameLogic_io_spriteYPosition_59; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_60 = gameLogic_io_spriteYPosition_60; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_61 = gameLogic_io_spriteYPosition_61; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_62 = gameLogic_io_spriteYPosition_62; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteYPosition_63 = gameLogic_io_spriteYPosition_63; // @[\\src\\main\\scala\\GameTop.scala 126:39]
  assign graphicEngineVGA_io_spriteVisible_3 = gameLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_4 = gameLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_5 = gameLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_6 = gameLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_7 = gameLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_8 = gameLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_9 = gameLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_10 = gameLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_11 = gameLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_12 = gameLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_13 = gameLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_14 = gameLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_15 = gameLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_16 = gameLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_17 = gameLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_18 = gameLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_19 = gameLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_20 = gameLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_21 = gameLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_22 = gameLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_23 = gameLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_24 = gameLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_25 = gameLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_26 = gameLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_27 = gameLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_28 = gameLogic_io_spriteVisible_28; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_29 = gameLogic_io_spriteVisible_29; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_30 = gameLogic_io_spriteVisible_30; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_31 = gameLogic_io_spriteVisible_31; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_32 = gameLogic_io_spriteVisible_32; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_33 = gameLogic_io_spriteVisible_33; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_34 = gameLogic_io_spriteVisible_34; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_35 = gameLogic_io_spriteVisible_35; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_36 = gameLogic_io_spriteVisible_36; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_37 = gameLogic_io_spriteVisible_37; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_38 = gameLogic_io_spriteVisible_38; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_39 = gameLogic_io_spriteVisible_39; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_40 = gameLogic_io_spriteVisible_40; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_41 = gameLogic_io_spriteVisible_41; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_42 = gameLogic_io_spriteVisible_42; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_43 = gameLogic_io_spriteVisible_43; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_44 = gameLogic_io_spriteVisible_44; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_45 = gameLogic_io_spriteVisible_45; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_46 = gameLogic_io_spriteVisible_46; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_47 = gameLogic_io_spriteVisible_47; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_48 = gameLogic_io_spriteVisible_48; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_49 = gameLogic_io_spriteVisible_49; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_50 = gameLogic_io_spriteVisible_50; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_51 = gameLogic_io_spriteVisible_51; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_52 = gameLogic_io_spriteVisible_52; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_53 = gameLogic_io_spriteVisible_53; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_54 = gameLogic_io_spriteVisible_54; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_55 = gameLogic_io_spriteVisible_55; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_56 = gameLogic_io_spriteVisible_56; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_57 = gameLogic_io_spriteVisible_57; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_58 = gameLogic_io_spriteVisible_58; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_59 = gameLogic_io_spriteVisible_59; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_60 = gameLogic_io_spriteVisible_60; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_61 = gameLogic_io_spriteVisible_61; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_62 = gameLogic_io_spriteVisible_62; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteVisible_63 = gameLogic_io_spriteVisible_63; // @[\\src\\main\\scala\\GameTop.scala 127:37]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_16 = gameLogic_io_spriteScaleUpHorizontal_16; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_17 = gameLogic_io_spriteScaleUpHorizontal_17; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_18 = gameLogic_io_spriteScaleUpHorizontal_18; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_19 = gameLogic_io_spriteScaleUpHorizontal_19; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_20 = gameLogic_io_spriteScaleUpHorizontal_20; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_21 = gameLogic_io_spriteScaleUpHorizontal_21; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_22 = gameLogic_io_spriteScaleUpHorizontal_22; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_23 = gameLogic_io_spriteScaleUpHorizontal_23; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_24 = gameLogic_io_spriteScaleUpHorizontal_24; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_25 = gameLogic_io_spriteScaleUpHorizontal_25; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_26 = gameLogic_io_spriteScaleUpHorizontal_26; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_27 = gameLogic_io_spriteScaleUpHorizontal_27; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_28 = gameLogic_io_spriteScaleUpHorizontal_28; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_29 = gameLogic_io_spriteScaleUpHorizontal_29; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_30 = gameLogic_io_spriteScaleUpHorizontal_30; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_31 = gameLogic_io_spriteScaleUpHorizontal_31; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_32 = gameLogic_io_spriteScaleUpHorizontal_32; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_33 = gameLogic_io_spriteScaleUpHorizontal_33; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_34 = gameLogic_io_spriteScaleUpHorizontal_34; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_35 = gameLogic_io_spriteScaleUpHorizontal_35; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_36 = gameLogic_io_spriteScaleUpHorizontal_36; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_37 = gameLogic_io_spriteScaleUpHorizontal_37; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_38 = gameLogic_io_spriteScaleUpHorizontal_38; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_39 = gameLogic_io_spriteScaleUpHorizontal_39; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_40 = gameLogic_io_spriteScaleUpHorizontal_40; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_41 = gameLogic_io_spriteScaleUpHorizontal_41; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_42 = gameLogic_io_spriteScaleUpHorizontal_42; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_43 = gameLogic_io_spriteScaleUpHorizontal_43; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_44 = gameLogic_io_spriteScaleUpHorizontal_44; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_45 = gameLogic_io_spriteScaleUpHorizontal_45; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_58 = gameLogic_io_spriteScaleUpHorizontal_58; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_59 = gameLogic_io_spriteScaleUpHorizontal_59; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpHorizontal_60 = gameLogic_io_spriteScaleUpHorizontal_60; // @[\\src\\main\\scala\\GameTop.scala 132:47]
  assign graphicEngineVGA_io_spriteScaleUpVertical_16 = gameLogic_io_spriteScaleUpVertical_16; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_17 = gameLogic_io_spriteScaleUpVertical_17; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_18 = gameLogic_io_spriteScaleUpVertical_18; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_19 = gameLogic_io_spriteScaleUpVertical_19; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_20 = gameLogic_io_spriteScaleUpVertical_20; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_21 = gameLogic_io_spriteScaleUpVertical_21; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_22 = gameLogic_io_spriteScaleUpVertical_22; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_23 = gameLogic_io_spriteScaleUpVertical_23; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_24 = gameLogic_io_spriteScaleUpVertical_24; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_25 = gameLogic_io_spriteScaleUpVertical_25; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_26 = gameLogic_io_spriteScaleUpVertical_26; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_27 = gameLogic_io_spriteScaleUpVertical_27; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_28 = gameLogic_io_spriteScaleUpVertical_28; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_29 = gameLogic_io_spriteScaleUpVertical_29; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_30 = gameLogic_io_spriteScaleUpVertical_30; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_31 = gameLogic_io_spriteScaleUpVertical_31; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_32 = gameLogic_io_spriteScaleUpVertical_32; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_33 = gameLogic_io_spriteScaleUpVertical_33; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_34 = gameLogic_io_spriteScaleUpVertical_34; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_35 = gameLogic_io_spriteScaleUpVertical_35; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_36 = gameLogic_io_spriteScaleUpVertical_36; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_37 = gameLogic_io_spriteScaleUpVertical_37; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_38 = gameLogic_io_spriteScaleUpVertical_38; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_39 = gameLogic_io_spriteScaleUpVertical_39; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_40 = gameLogic_io_spriteScaleUpVertical_40; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_41 = gameLogic_io_spriteScaleUpVertical_41; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_42 = gameLogic_io_spriteScaleUpVertical_42; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_43 = gameLogic_io_spriteScaleUpVertical_43; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_44 = gameLogic_io_spriteScaleUpVertical_44; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_45 = gameLogic_io_spriteScaleUpVertical_45; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_58 = gameLogic_io_spriteScaleUpVertical_58; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_59 = gameLogic_io_spriteScaleUpVertical_59; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_spriteScaleUpVertical_60 = gameLogic_io_spriteScaleUpVertical_60; // @[\\src\\main\\scala\\GameTop.scala 134:45]
  assign graphicEngineVGA_io_viewBoxX = gameLogic_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 138:32]
  assign graphicEngineVGA_io_viewBoxY = gameLogic_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 139:32]
  assign graphicEngineVGA_io_frameUpdateDone = gameLogic_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 148:39]
  assign soundEngine_clock = clock;
  assign soundEngine_reset = reset;
  assign gameLogic_clock = clock;
  assign gameLogic_reset = resetReleaseCounter == 22'h3d08ff ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameTop.scala 83:67 84:18 86:18]
  assign gameLogic_io_btnC = btnCState; // @[\\src\\main\\scala\\GameTop.scala 98:21]
  assign gameLogic_io_btnU = btnUState; // @[\\src\\main\\scala\\GameTop.scala 99:21]
  assign gameLogic_io_btnL = btnLState; // @[\\src\\main\\scala\\GameTop.scala 100:21]
  assign gameLogic_io_btnR = btnRState; // @[\\src\\main\\scala\\GameTop.scala 101:21]
  assign gameLogic_io_btnD = btnDState; // @[\\src\\main\\scala\\GameTop.scala 102:21]
  assign gameLogic_io_newFrame = graphicEngineVGA_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 147:25]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 68:32]
      debounceCounter <= 21'h0; // @[\\src\\main\\scala\\GameTop.scala 68:32]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 70:57]
      debounceCounter <= 21'h0; // @[\\src\\main\\scala\\GameTop.scala 71:21]
    end else begin
      debounceCounter <= _debounceCounter_T_1; // @[\\src\\main\\scala\\GameTop.scala 74:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 81:36]
      resetReleaseCounter <= 22'h0; // @[\\src\\main\\scala\\GameTop.scala 81:36]
    end else if (!(resetReleaseCounter == 22'h3d08ff)) begin // @[\\src\\main\\scala\\GameTop.scala 83:67]
      resetReleaseCounter <= _resetReleaseCounter_T_1; // @[\\src\\main\\scala\\GameTop.scala 87:25]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnCState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnCState_pipeReg_0 <= btnCState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnCState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnCState_pipeReg_1 <= btnCState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnCState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnCState_pipeReg_2 <= io_btnC; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 93:28]
      btnCState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 93:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 93:28]
      btnCState <= btnCState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 93:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_0 <= btnUState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_1 <= btnUState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_2 <= io_btnU; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 94:28]
      btnUState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 94:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 94:28]
      btnUState <= btnUState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 94:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_0 <= btnLState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_1 <= btnLState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_2 <= io_btnL; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 95:28]
      btnLState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 95:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 95:28]
      btnLState <= btnLState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 95:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_0 <= btnRState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_1 <= btnRState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_2 <= io_btnR; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 96:28]
      btnRState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 96:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 96:28]
      btnRState <= btnRState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 96:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_0 <= btnDState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_1 <= btnDState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_2 <= io_btnD; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 97:28]
      btnDState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 97:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 97:28]
      btnDState <= btnDState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 97:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounceCounter = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  resetReleaseCounter = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btnCState_pipeReg_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  btnCState_pipeReg_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  btnCState_pipeReg_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  btnCState = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  btnUState_pipeReg_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  btnUState_pipeReg_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  btnUState_pipeReg_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btnUState = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  btnLState_pipeReg_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  btnLState_pipeReg_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  btnLState_pipeReg_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btnLState = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  btnRState_pipeReg_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  btnRState_pipeReg_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  btnRState_pipeReg_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  btnRState = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  btnDState_pipeReg_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  btnDState_pipeReg_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  btnDState_pipeReg_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  btnDState = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input        clock,
  input        reset,
  input        io_btnC, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnU, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnL, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnR, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnD, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaRed, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaGreen, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaBlue, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_Hsync, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_Vsync, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_0, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_1, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_2, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_3, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_4, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_5, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_6, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_7, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_0, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_1, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_2, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_3, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_4, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_5, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_6, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_7, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_missingFrameError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_backBufferWriteError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_viewBoxOutOfRangeError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_soundOut // @[\\src\\main\\scala\\Top.scala 14:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  gameTop_clock; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_reset; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnC; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnU; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnL; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnR; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnD; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaRed; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaBlue; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaGreen; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_Hsync; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_Vsync; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_missingFrameError; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\Top.scala 44:23]
  reg  syncResetInput_REG; // @[\\src\\main\\scala\\Top.scala 49:48]
  reg  syncResetInput_REG_1; // @[\\src\\main\\scala\\Top.scala 49:40]
  reg  syncResetInput_REG_2; // @[\\src\\main\\scala\\Top.scala 49:32]
  reg  pipeResetReg_0; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_1; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_2; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_3; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_4; // @[\\src\\main\\scala\\Top.scala 54:25]
  wire [4:0] _gameTop_reset_T = {pipeResetReg_4,pipeResetReg_3,pipeResetReg_2,pipeResetReg_1,pipeResetReg_0}; // @[\\src\\main\\scala\\Top.scala 59:33]
  GameTop gameTop ( // @[\\src\\main\\scala\\Top.scala 44:23]
    .clock(gameTop_clock),
    .reset(gameTop_reset),
    .io_btnC(gameTop_io_btnC),
    .io_btnU(gameTop_io_btnU),
    .io_btnL(gameTop_io_btnL),
    .io_btnR(gameTop_io_btnR),
    .io_btnD(gameTop_io_btnD),
    .io_vgaRed(gameTop_io_vgaRed),
    .io_vgaBlue(gameTop_io_vgaBlue),
    .io_vgaGreen(gameTop_io_vgaGreen),
    .io_Hsync(gameTop_io_Hsync),
    .io_Vsync(gameTop_io_Vsync),
    .io_missingFrameError(gameTop_io_missingFrameError),
    .io_viewBoxOutOfRangeError(gameTop_io_viewBoxOutOfRangeError)
  );
  assign io_vgaRed = gameTop_io_vgaRed; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_vgaGreen = gameTop_io_vgaGreen; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_vgaBlue = gameTop_io_vgaBlue; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_Hsync = gameTop_io_Hsync; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_Vsync = gameTop_io_Vsync; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_0 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_1 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_2 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_3 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_4 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_5 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_6 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_7 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_missingFrameError = gameTop_io_missingFrameError; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_backBufferWriteError = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_viewBoxOutOfRangeError = gameTop_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_soundOut = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_clock = clock;
  assign gameTop_reset = |_gameTop_reset_T; // @[\\src\\main\\scala\\Top.scala 59:40]
  assign gameTop_io_btnC = io_btnC; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnU = io_btnU; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnL = io_btnL; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnR = io_btnR; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnD = io_btnD; // @[\\src\\main\\scala\\Top.scala 62:14]
  always @(posedge clock) begin
    syncResetInput_REG <= reset; // @[\\src\\main\\scala\\Top.scala 49:48]
    syncResetInput_REG_1 <= syncResetInput_REG; // @[\\src\\main\\scala\\Top.scala 49:40]
    syncResetInput_REG_2 <= syncResetInput_REG_1; // @[\\src\\main\\scala\\Top.scala 49:32]
    pipeResetReg_0 <= pipeResetReg_1; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_1 <= pipeResetReg_2; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_2 <= pipeResetReg_3; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_3 <= pipeResetReg_4; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_4 <= ~syncResetInput_REG_2; // @[\\src\\main\\scala\\Top.scala 49:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  syncResetInput_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  syncResetInput_REG_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  syncResetInput_REG_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pipeResetReg_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pipeResetReg_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pipeResetReg_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pipeResetReg_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pipeResetReg_4 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
